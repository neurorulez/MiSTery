
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"00",x"60"),
     1 => (x"08",x"08",x"08",x"00"),
     2 => (x"00",x"08",x"08",x"08"),
     3 => (x"60",x"00",x"00",x"00"),
     4 => (x"00",x"00",x"00",x"60"),
     5 => (x"18",x"30",x"60",x"40"),
     6 => (x"01",x"03",x"06",x"0c"),
     7 => (x"59",x"7f",x"3e",x"00"),
     8 => (x"00",x"3e",x"7f",x"4d"),
     9 => (x"7f",x"06",x"04",x"00"),
    10 => (x"00",x"00",x"00",x"7f"),
    11 => (x"71",x"63",x"42",x"00"),
    12 => (x"00",x"46",x"4f",x"59"),
    13 => (x"49",x"63",x"22",x"00"),
    14 => (x"00",x"36",x"7f",x"49"),
    15 => (x"13",x"16",x"1c",x"18"),
    16 => (x"00",x"10",x"7f",x"7f"),
    17 => (x"45",x"67",x"27",x"00"),
    18 => (x"00",x"39",x"7d",x"45"),
    19 => (x"4b",x"7e",x"3c",x"00"),
    20 => (x"00",x"30",x"79",x"49"),
    21 => (x"71",x"01",x"01",x"00"),
    22 => (x"00",x"07",x"0f",x"79"),
    23 => (x"49",x"7f",x"36",x"00"),
    24 => (x"00",x"36",x"7f",x"49"),
    25 => (x"49",x"4f",x"06",x"00"),
    26 => (x"00",x"1e",x"3f",x"69"),
    27 => (x"66",x"00",x"00",x"00"),
    28 => (x"00",x"00",x"00",x"66"),
    29 => (x"e6",x"80",x"00",x"00"),
    30 => (x"00",x"00",x"00",x"66"),
    31 => (x"14",x"08",x"08",x"00"),
    32 => (x"00",x"22",x"22",x"14"),
    33 => (x"14",x"14",x"14",x"00"),
    34 => (x"00",x"14",x"14",x"14"),
    35 => (x"14",x"22",x"22",x"00"),
    36 => (x"00",x"08",x"08",x"14"),
    37 => (x"51",x"03",x"02",x"00"),
    38 => (x"00",x"06",x"0f",x"59"),
    39 => (x"5d",x"41",x"7f",x"3e"),
    40 => (x"00",x"1e",x"1f",x"55"),
    41 => (x"09",x"7f",x"7e",x"00"),
    42 => (x"00",x"7e",x"7f",x"09"),
    43 => (x"49",x"7f",x"7f",x"00"),
    44 => (x"00",x"36",x"7f",x"49"),
    45 => (x"63",x"3e",x"1c",x"00"),
    46 => (x"00",x"41",x"41",x"41"),
    47 => (x"41",x"7f",x"7f",x"00"),
    48 => (x"00",x"1c",x"3e",x"63"),
    49 => (x"49",x"7f",x"7f",x"00"),
    50 => (x"00",x"41",x"41",x"49"),
    51 => (x"09",x"7f",x"7f",x"00"),
    52 => (x"00",x"01",x"01",x"09"),
    53 => (x"41",x"7f",x"3e",x"00"),
    54 => (x"00",x"7a",x"7b",x"49"),
    55 => (x"08",x"7f",x"7f",x"00"),
    56 => (x"00",x"7f",x"7f",x"08"),
    57 => (x"7f",x"41",x"00",x"00"),
    58 => (x"00",x"00",x"41",x"7f"),
    59 => (x"40",x"60",x"20",x"00"),
    60 => (x"00",x"3f",x"7f",x"40"),
    61 => (x"1c",x"08",x"7f",x"7f"),
    62 => (x"00",x"41",x"63",x"36"),
    63 => (x"40",x"7f",x"7f",x"00"),
    64 => (x"00",x"40",x"40",x"40"),
    65 => (x"0c",x"06",x"7f",x"7f"),
    66 => (x"00",x"7f",x"7f",x"06"),
    67 => (x"0c",x"06",x"7f",x"7f"),
    68 => (x"00",x"7f",x"7f",x"18"),
    69 => (x"41",x"7f",x"3e",x"00"),
    70 => (x"00",x"3e",x"7f",x"41"),
    71 => (x"09",x"7f",x"7f",x"00"),
    72 => (x"00",x"06",x"0f",x"09"),
    73 => (x"61",x"41",x"7f",x"3e"),
    74 => (x"00",x"40",x"7e",x"7f"),
    75 => (x"09",x"7f",x"7f",x"00"),
    76 => (x"00",x"66",x"7f",x"19"),
    77 => (x"4d",x"6f",x"26",x"00"),
    78 => (x"00",x"32",x"7b",x"59"),
    79 => (x"7f",x"01",x"01",x"00"),
    80 => (x"00",x"01",x"01",x"7f"),
    81 => (x"40",x"7f",x"3f",x"00"),
    82 => (x"00",x"3f",x"7f",x"40"),
    83 => (x"70",x"3f",x"0f",x"00"),
    84 => (x"00",x"0f",x"3f",x"70"),
    85 => (x"18",x"30",x"7f",x"7f"),
    86 => (x"00",x"7f",x"7f",x"30"),
    87 => (x"1c",x"36",x"63",x"41"),
    88 => (x"41",x"63",x"36",x"1c"),
    89 => (x"7c",x"06",x"03",x"01"),
    90 => (x"01",x"03",x"06",x"7c"),
    91 => (x"4d",x"59",x"71",x"61"),
    92 => (x"00",x"41",x"43",x"47"),
    93 => (x"7f",x"7f",x"00",x"00"),
    94 => (x"00",x"00",x"41",x"41"),
    95 => (x"0c",x"06",x"03",x"01"),
    96 => (x"40",x"60",x"30",x"18"),
    97 => (x"41",x"41",x"00",x"00"),
    98 => (x"00",x"00",x"7f",x"7f"),
    99 => (x"03",x"06",x"0c",x"08"),
   100 => (x"00",x"08",x"0c",x"06"),
   101 => (x"80",x"80",x"80",x"80"),
   102 => (x"00",x"80",x"80",x"80"),
   103 => (x"03",x"00",x"00",x"00"),
   104 => (x"00",x"00",x"04",x"07"),
   105 => (x"54",x"74",x"20",x"00"),
   106 => (x"00",x"78",x"7c",x"54"),
   107 => (x"44",x"7f",x"7f",x"00"),
   108 => (x"00",x"38",x"7c",x"44"),
   109 => (x"44",x"7c",x"38",x"00"),
   110 => (x"00",x"00",x"44",x"44"),
   111 => (x"44",x"7c",x"38",x"00"),
   112 => (x"00",x"7f",x"7f",x"44"),
   113 => (x"54",x"7c",x"38",x"00"),
   114 => (x"00",x"18",x"5c",x"54"),
   115 => (x"7f",x"7e",x"04",x"00"),
   116 => (x"00",x"00",x"05",x"05"),
   117 => (x"a4",x"bc",x"18",x"00"),
   118 => (x"00",x"7c",x"fc",x"a4"),
   119 => (x"04",x"7f",x"7f",x"00"),
   120 => (x"00",x"78",x"7c",x"04"),
   121 => (x"3d",x"00",x"00",x"00"),
   122 => (x"00",x"00",x"40",x"7d"),
   123 => (x"80",x"80",x"80",x"00"),
   124 => (x"00",x"00",x"7d",x"fd"),
   125 => (x"10",x"7f",x"7f",x"00"),
   126 => (x"00",x"44",x"6c",x"38"),
   127 => (x"3f",x"00",x"00",x"00"),
   128 => (x"00",x"00",x"40",x"7f"),
   129 => (x"18",x"0c",x"7c",x"7c"),
   130 => (x"00",x"78",x"7c",x"0c"),
   131 => (x"04",x"7c",x"7c",x"00"),
   132 => (x"00",x"78",x"7c",x"04"),
   133 => (x"44",x"7c",x"38",x"00"),
   134 => (x"00",x"38",x"7c",x"44"),
   135 => (x"24",x"fc",x"fc",x"00"),
   136 => (x"00",x"18",x"3c",x"24"),
   137 => (x"24",x"3c",x"18",x"00"),
   138 => (x"00",x"fc",x"fc",x"24"),
   139 => (x"04",x"7c",x"7c",x"00"),
   140 => (x"00",x"08",x"0c",x"04"),
   141 => (x"54",x"5c",x"48",x"00"),
   142 => (x"00",x"20",x"74",x"54"),
   143 => (x"7f",x"3f",x"04",x"00"),
   144 => (x"00",x"00",x"44",x"44"),
   145 => (x"40",x"7c",x"3c",x"00"),
   146 => (x"00",x"7c",x"7c",x"40"),
   147 => (x"60",x"3c",x"1c",x"00"),
   148 => (x"00",x"1c",x"3c",x"60"),
   149 => (x"30",x"60",x"7c",x"3c"),
   150 => (x"00",x"3c",x"7c",x"60"),
   151 => (x"10",x"38",x"6c",x"44"),
   152 => (x"00",x"44",x"6c",x"38"),
   153 => (x"e0",x"bc",x"1c",x"00"),
   154 => (x"00",x"1c",x"3c",x"60"),
   155 => (x"74",x"64",x"44",x"00"),
   156 => (x"00",x"44",x"4c",x"5c"),
   157 => (x"3e",x"08",x"08",x"00"),
   158 => (x"00",x"41",x"41",x"77"),
   159 => (x"7f",x"00",x"00",x"00"),
   160 => (x"00",x"00",x"00",x"7f"),
   161 => (x"77",x"41",x"41",x"00"),
   162 => (x"00",x"08",x"08",x"3e"),
   163 => (x"03",x"01",x"01",x"02"),
   164 => (x"00",x"01",x"02",x"02"),
   165 => (x"7f",x"7f",x"7f",x"7f"),
   166 => (x"00",x"7f",x"7f",x"7f"),
   167 => (x"1c",x"1c",x"08",x"08"),
   168 => (x"7f",x"7f",x"3e",x"3e"),
   169 => (x"3e",x"3e",x"7f",x"7f"),
   170 => (x"08",x"08",x"1c",x"1c"),
   171 => (x"7c",x"18",x"10",x"00"),
   172 => (x"00",x"10",x"18",x"7c"),
   173 => (x"7c",x"30",x"10",x"00"),
   174 => (x"00",x"10",x"30",x"7c"),
   175 => (x"60",x"60",x"30",x"10"),
   176 => (x"00",x"06",x"1e",x"78"),
   177 => (x"18",x"3c",x"66",x"42"),
   178 => (x"00",x"42",x"66",x"3c"),
   179 => (x"c2",x"6a",x"38",x"78"),
   180 => (x"00",x"38",x"6c",x"c6"),
   181 => (x"60",x"00",x"00",x"60"),
   182 => (x"00",x"60",x"00",x"00"),
   183 => (x"5c",x"5b",x"5e",x"0e"),
   184 => (x"86",x"fc",x"0e",x"5d"),
   185 => (x"ca",x"c3",x"7e",x"71"),
   186 => (x"c0",x"4c",x"bf",x"c0"),
   187 => (x"c4",x"1e",x"c0",x"4b"),
   188 => (x"c4",x"02",x"ab",x"66"),
   189 => (x"c2",x"4d",x"c0",x"87"),
   190 => (x"75",x"4d",x"c1",x"87"),
   191 => (x"ee",x"49",x"73",x"1e"),
   192 => (x"86",x"c8",x"87",x"e3"),
   193 => (x"ef",x"49",x"e0",x"c0"),
   194 => (x"a4",x"c4",x"87",x"ec"),
   195 => (x"f0",x"49",x"6a",x"4a"),
   196 => (x"ca",x"f1",x"87",x"f3"),
   197 => (x"c1",x"84",x"cc",x"87"),
   198 => (x"ab",x"b7",x"c8",x"83"),
   199 => (x"87",x"cd",x"ff",x"04"),
   200 => (x"4d",x"26",x"8e",x"fc"),
   201 => (x"4b",x"26",x"4c",x"26"),
   202 => (x"71",x"1e",x"4f",x"26"),
   203 => (x"c4",x"ca",x"c3",x"4a"),
   204 => (x"c4",x"ca",x"c3",x"5a"),
   205 => (x"49",x"78",x"c7",x"48"),
   206 => (x"26",x"87",x"e1",x"fe"),
   207 => (x"1e",x"73",x"1e",x"4f"),
   208 => (x"0b",x"fc",x"4b",x"71"),
   209 => (x"4a",x"73",x"0b",x"7b"),
   210 => (x"c0",x"c1",x"9a",x"c1"),
   211 => (x"c7",x"ed",x"49",x"a2"),
   212 => (x"d0",x"da",x"c2",x"87"),
   213 => (x"26",x"4b",x"26",x"5b"),
   214 => (x"4a",x"71",x"1e",x"4f"),
   215 => (x"72",x"1e",x"66",x"c4"),
   216 => (x"87",x"fb",x"eb",x"49"),
   217 => (x"4f",x"26",x"8e",x"fc"),
   218 => (x"48",x"d4",x"ff",x"1e"),
   219 => (x"ff",x"78",x"ff",x"c3"),
   220 => (x"e1",x"c0",x"48",x"d0"),
   221 => (x"48",x"d4",x"ff",x"78"),
   222 => (x"48",x"71",x"78",x"c1"),
   223 => (x"d4",x"ff",x"30",x"c4"),
   224 => (x"d0",x"ff",x"78",x"08"),
   225 => (x"78",x"e0",x"c0",x"48"),
   226 => (x"5e",x"0e",x"4f",x"26"),
   227 => (x"0e",x"5d",x"5c",x"5b"),
   228 => (x"7e",x"c0",x"86",x"f4"),
   229 => (x"ec",x"48",x"a6",x"c8"),
   230 => (x"80",x"fc",x"78",x"bf"),
   231 => (x"bf",x"c0",x"ca",x"c3"),
   232 => (x"c8",x"ca",x"c3",x"78"),
   233 => (x"bf",x"e8",x"4c",x"bf"),
   234 => (x"cc",x"da",x"c2",x"4d"),
   235 => (x"ef",x"e4",x"49",x"bf"),
   236 => (x"e8",x"49",x"c7",x"87"),
   237 => (x"49",x"70",x"87",x"f1"),
   238 => (x"d0",x"05",x"99",x"c2"),
   239 => (x"c4",x"da",x"c2",x"87"),
   240 => (x"b9",x"ff",x"49",x"bf"),
   241 => (x"c1",x"99",x"66",x"c8"),
   242 => (x"f9",x"c1",x"02",x"99"),
   243 => (x"49",x"e8",x"cf",x"87"),
   244 => (x"70",x"87",x"fd",x"ca"),
   245 => (x"e8",x"49",x"c7",x"4b"),
   246 => (x"98",x"70",x"87",x"cd"),
   247 => (x"c8",x"87",x"c9",x"05"),
   248 => (x"99",x"c1",x"49",x"66"),
   249 => (x"87",x"fe",x"c0",x"02"),
   250 => (x"ec",x"48",x"a6",x"c8"),
   251 => (x"ef",x"e3",x"78",x"bf"),
   252 => (x"ca",x"49",x"73",x"87"),
   253 => (x"98",x"70",x"87",x"e6"),
   254 => (x"c2",x"87",x"d7",x"02"),
   255 => (x"49",x"bf",x"c0",x"da"),
   256 => (x"da",x"c2",x"b9",x"c1"),
   257 => (x"fd",x"71",x"59",x"c4"),
   258 => (x"e8",x"cf",x"87",x"de"),
   259 => (x"87",x"c0",x"ca",x"49"),
   260 => (x"49",x"c7",x"4b",x"70"),
   261 => (x"70",x"87",x"d0",x"e7"),
   262 => (x"cb",x"ff",x"05",x"98"),
   263 => (x"49",x"66",x"c8",x"87"),
   264 => (x"ff",x"05",x"99",x"c1"),
   265 => (x"da",x"c2",x"87",x"c2"),
   266 => (x"c1",x"4a",x"bf",x"cc"),
   267 => (x"d0",x"da",x"c2",x"ba"),
   268 => (x"7a",x"0a",x"fc",x"5a"),
   269 => (x"c1",x"9a",x"c1",x"0a"),
   270 => (x"e9",x"49",x"a2",x"c0"),
   271 => (x"da",x"c1",x"87",x"da"),
   272 => (x"87",x"e3",x"e6",x"49"),
   273 => (x"da",x"c2",x"7e",x"c1"),
   274 => (x"66",x"c8",x"48",x"c4"),
   275 => (x"cc",x"da",x"c2",x"78"),
   276 => (x"e9",x"c0",x"05",x"bf"),
   277 => (x"c3",x"49",x"75",x"87"),
   278 => (x"1e",x"71",x"99",x"ff"),
   279 => (x"f8",x"fb",x"49",x"c0"),
   280 => (x"c8",x"49",x"75",x"87"),
   281 => (x"1e",x"71",x"29",x"b7"),
   282 => (x"ec",x"fb",x"49",x"c1"),
   283 => (x"c3",x"86",x"c8",x"87"),
   284 => (x"f2",x"e5",x"49",x"fd"),
   285 => (x"49",x"fa",x"c3",x"87"),
   286 => (x"c7",x"87",x"ec",x"e5"),
   287 => (x"49",x"75",x"87",x"f4"),
   288 => (x"c8",x"99",x"ff",x"c3"),
   289 => (x"b5",x"71",x"2d",x"b7"),
   290 => (x"c0",x"02",x"9d",x"75"),
   291 => (x"a6",x"c8",x"87",x"e4"),
   292 => (x"bf",x"c8",x"ff",x"48"),
   293 => (x"49",x"66",x"c8",x"78"),
   294 => (x"bf",x"c8",x"da",x"c2"),
   295 => (x"a9",x"e0",x"c2",x"89"),
   296 => (x"87",x"c4",x"c0",x"03"),
   297 => (x"87",x"d0",x"4d",x"c0"),
   298 => (x"48",x"c8",x"da",x"c2"),
   299 => (x"c0",x"78",x"66",x"c8"),
   300 => (x"da",x"c2",x"87",x"c6"),
   301 => (x"78",x"c0",x"48",x"c8"),
   302 => (x"99",x"c8",x"49",x"75"),
   303 => (x"87",x"ce",x"c0",x"05"),
   304 => (x"e4",x"49",x"f5",x"c3"),
   305 => (x"49",x"70",x"87",x"e1"),
   306 => (x"c0",x"02",x"99",x"c2"),
   307 => (x"ca",x"c3",x"87",x"e7"),
   308 => (x"c0",x"02",x"bf",x"c4"),
   309 => (x"c1",x"48",x"87",x"ca"),
   310 => (x"c8",x"ca",x"c3",x"88"),
   311 => (x"87",x"d3",x"c0",x"58"),
   312 => (x"c1",x"48",x"66",x"c4"),
   313 => (x"7e",x"70",x"80",x"e0"),
   314 => (x"c0",x"02",x"bf",x"6e"),
   315 => (x"ff",x"4b",x"87",x"c5"),
   316 => (x"c1",x"0f",x"73",x"49"),
   317 => (x"c4",x"49",x"75",x"7e"),
   318 => (x"ce",x"c0",x"05",x"99"),
   319 => (x"49",x"f2",x"c3",x"87"),
   320 => (x"70",x"87",x"e4",x"e3"),
   321 => (x"02",x"99",x"c2",x"49"),
   322 => (x"c3",x"87",x"ea",x"c0"),
   323 => (x"7e",x"bf",x"c4",x"ca"),
   324 => (x"a8",x"b7",x"c7",x"48"),
   325 => (x"87",x"cb",x"c0",x"03"),
   326 => (x"80",x"c1",x"48",x"6e"),
   327 => (x"58",x"c8",x"ca",x"c3"),
   328 => (x"c4",x"87",x"d0",x"c0"),
   329 => (x"e0",x"c1",x"4a",x"66"),
   330 => (x"c0",x"02",x"6a",x"82"),
   331 => (x"fe",x"4b",x"87",x"c5"),
   332 => (x"c1",x"0f",x"73",x"49"),
   333 => (x"49",x"fd",x"c3",x"7e"),
   334 => (x"70",x"87",x"ec",x"e2"),
   335 => (x"02",x"99",x"c2",x"49"),
   336 => (x"c3",x"87",x"e6",x"c0"),
   337 => (x"02",x"bf",x"c4",x"ca"),
   338 => (x"c3",x"87",x"c9",x"c0"),
   339 => (x"c0",x"48",x"c4",x"ca"),
   340 => (x"87",x"d3",x"c0",x"78"),
   341 => (x"c1",x"48",x"66",x"c4"),
   342 => (x"7e",x"70",x"80",x"e0"),
   343 => (x"c0",x"02",x"bf",x"6e"),
   344 => (x"fd",x"4b",x"87",x"c5"),
   345 => (x"c1",x"0f",x"73",x"49"),
   346 => (x"49",x"fa",x"c3",x"7e"),
   347 => (x"70",x"87",x"f8",x"e1"),
   348 => (x"02",x"99",x"c2",x"49"),
   349 => (x"c3",x"87",x"ea",x"c0"),
   350 => (x"48",x"bf",x"c4",x"ca"),
   351 => (x"03",x"a8",x"b7",x"c7"),
   352 => (x"c3",x"87",x"c9",x"c0"),
   353 => (x"c7",x"48",x"c4",x"ca"),
   354 => (x"87",x"d3",x"c0",x"78"),
   355 => (x"c1",x"48",x"66",x"c4"),
   356 => (x"7e",x"70",x"80",x"e0"),
   357 => (x"c0",x"02",x"bf",x"6e"),
   358 => (x"fc",x"4b",x"87",x"c5"),
   359 => (x"c1",x"0f",x"73",x"49"),
   360 => (x"c3",x"48",x"75",x"7e"),
   361 => (x"a6",x"cc",x"98",x"f0"),
   362 => (x"05",x"98",x"70",x"58"),
   363 => (x"c1",x"87",x"ce",x"c0"),
   364 => (x"f2",x"e0",x"49",x"da"),
   365 => (x"c2",x"49",x"70",x"87"),
   366 => (x"f9",x"c1",x"02",x"99"),
   367 => (x"49",x"e8",x"cf",x"87"),
   368 => (x"70",x"87",x"cd",x"c3"),
   369 => (x"fc",x"c9",x"c3",x"4b"),
   370 => (x"c3",x"50",x"c0",x"48"),
   371 => (x"bf",x"97",x"fc",x"c9"),
   372 => (x"87",x"d2",x"c1",x"05"),
   373 => (x"c0",x"05",x"66",x"c8"),
   374 => (x"da",x"c1",x"87",x"cc"),
   375 => (x"87",x"c7",x"e0",x"49"),
   376 => (x"c1",x"02",x"98",x"70"),
   377 => (x"bf",x"e8",x"87",x"c0"),
   378 => (x"ff",x"c3",x"49",x"4d"),
   379 => (x"2d",x"b7",x"c8",x"99"),
   380 => (x"db",x"ff",x"b5",x"71"),
   381 => (x"49",x"73",x"87",x"ea"),
   382 => (x"70",x"87",x"e1",x"c2"),
   383 => (x"c6",x"c0",x"02",x"98"),
   384 => (x"fc",x"c9",x"c3",x"87"),
   385 => (x"c3",x"50",x"c1",x"48"),
   386 => (x"bf",x"97",x"fc",x"c9"),
   387 => (x"87",x"d6",x"c0",x"05"),
   388 => (x"f0",x"c3",x"49",x"75"),
   389 => (x"cd",x"ff",x"05",x"99"),
   390 => (x"49",x"da",x"c1",x"87"),
   391 => (x"87",x"c7",x"df",x"ff"),
   392 => (x"ff",x"05",x"98",x"70"),
   393 => (x"ca",x"c3",x"87",x"c0"),
   394 => (x"4b",x"49",x"bf",x"c4"),
   395 => (x"66",x"c4",x"93",x"cc"),
   396 => (x"71",x"4b",x"6b",x"83"),
   397 => (x"9c",x"74",x"0f",x"73"),
   398 => (x"87",x"e9",x"c0",x"02"),
   399 => (x"e4",x"c0",x"02",x"6c"),
   400 => (x"ff",x"49",x"6c",x"87"),
   401 => (x"70",x"87",x"e0",x"de"),
   402 => (x"02",x"99",x"c1",x"49"),
   403 => (x"c4",x"87",x"cb",x"c0"),
   404 => (x"ca",x"c3",x"4b",x"a4"),
   405 => (x"6b",x"49",x"bf",x"c4"),
   406 => (x"84",x"c8",x"0f",x"4b"),
   407 => (x"87",x"c5",x"c0",x"02"),
   408 => (x"dc",x"ff",x"05",x"6c"),
   409 => (x"c0",x"02",x"6e",x"87"),
   410 => (x"ca",x"c3",x"87",x"c8"),
   411 => (x"f1",x"49",x"bf",x"c4"),
   412 => (x"8e",x"f4",x"87",x"ea"),
   413 => (x"4c",x"26",x"4d",x"26"),
   414 => (x"4f",x"26",x"4b",x"26"),
   415 => (x"00",x"00",x"00",x"10"),
   416 => (x"00",x"00",x"00",x"00"),
   417 => (x"00",x"00",x"00",x"00"),
   418 => (x"00",x"00",x"00",x"00"),
   419 => (x"00",x"00",x"00",x"00"),
   420 => (x"ff",x"4a",x"71",x"1e"),
   421 => (x"72",x"49",x"bf",x"c8"),
   422 => (x"4f",x"26",x"48",x"a1"),
   423 => (x"bf",x"c8",x"ff",x"1e"),
   424 => (x"c0",x"c0",x"fe",x"89"),
   425 => (x"a9",x"c0",x"c0",x"c0"),
   426 => (x"c0",x"87",x"c4",x"01"),
   427 => (x"c1",x"87",x"c2",x"4a"),
   428 => (x"26",x"48",x"72",x"4a"),
   429 => (x"5b",x"5e",x"0e",x"4f"),
   430 => (x"71",x"0e",x"5d",x"5c"),
   431 => (x"4c",x"d4",x"ff",x"4b"),
   432 => (x"c0",x"48",x"66",x"d0"),
   433 => (x"ff",x"49",x"d6",x"78"),
   434 => (x"c3",x"87",x"d9",x"dd"),
   435 => (x"49",x"6c",x"7c",x"ff"),
   436 => (x"71",x"99",x"ff",x"c3"),
   437 => (x"f0",x"c3",x"49",x"4d"),
   438 => (x"a9",x"e0",x"c1",x"99"),
   439 => (x"c3",x"87",x"cb",x"05"),
   440 => (x"48",x"6c",x"7c",x"ff"),
   441 => (x"66",x"d0",x"98",x"c3"),
   442 => (x"ff",x"c3",x"78",x"08"),
   443 => (x"49",x"4a",x"6c",x"7c"),
   444 => (x"ff",x"c3",x"31",x"c8"),
   445 => (x"71",x"4a",x"6c",x"7c"),
   446 => (x"c8",x"49",x"72",x"b2"),
   447 => (x"7c",x"ff",x"c3",x"31"),
   448 => (x"b2",x"71",x"4a",x"6c"),
   449 => (x"31",x"c8",x"49",x"72"),
   450 => (x"6c",x"7c",x"ff",x"c3"),
   451 => (x"ff",x"b2",x"71",x"4a"),
   452 => (x"e0",x"c0",x"48",x"d0"),
   453 => (x"02",x"9b",x"73",x"78"),
   454 => (x"7b",x"72",x"87",x"c2"),
   455 => (x"4d",x"26",x"48",x"75"),
   456 => (x"4b",x"26",x"4c",x"26"),
   457 => (x"26",x"1e",x"4f",x"26"),
   458 => (x"5b",x"5e",x"0e",x"4f"),
   459 => (x"86",x"f8",x"0e",x"5c"),
   460 => (x"a6",x"c8",x"1e",x"76"),
   461 => (x"87",x"fd",x"fd",x"49"),
   462 => (x"4b",x"70",x"86",x"c4"),
   463 => (x"a8",x"c2",x"48",x"6e"),
   464 => (x"87",x"fb",x"c2",x"03"),
   465 => (x"f0",x"c3",x"4a",x"73"),
   466 => (x"aa",x"d0",x"c1",x"9a"),
   467 => (x"c1",x"87",x"c7",x"02"),
   468 => (x"c2",x"05",x"aa",x"e0"),
   469 => (x"49",x"73",x"87",x"e9"),
   470 => (x"c3",x"02",x"99",x"c8"),
   471 => (x"87",x"c6",x"ff",x"87"),
   472 => (x"9c",x"c3",x"4c",x"73"),
   473 => (x"c1",x"05",x"ac",x"c2"),
   474 => (x"66",x"c4",x"87",x"c4"),
   475 => (x"71",x"31",x"c9",x"49"),
   476 => (x"4a",x"66",x"c4",x"1e"),
   477 => (x"c3",x"92",x"cc",x"c1"),
   478 => (x"72",x"49",x"cc",x"ca"),
   479 => (x"cb",x"cd",x"fe",x"81"),
   480 => (x"ff",x"49",x"d8",x"87"),
   481 => (x"c8",x"87",x"dd",x"da"),
   482 => (x"f6",x"c2",x"1e",x"c0"),
   483 => (x"e6",x"fd",x"49",x"e8"),
   484 => (x"d0",x"ff",x"87",x"e1"),
   485 => (x"78",x"e0",x"c0",x"48"),
   486 => (x"1e",x"e8",x"f6",x"c2"),
   487 => (x"c1",x"4a",x"66",x"cc"),
   488 => (x"ca",x"c3",x"92",x"cc"),
   489 => (x"81",x"72",x"49",x"cc"),
   490 => (x"87",x"e1",x"cb",x"fe"),
   491 => (x"ac",x"c1",x"86",x"cc"),
   492 => (x"87",x"cb",x"c1",x"05"),
   493 => (x"fd",x"49",x"ee",x"c0"),
   494 => (x"c4",x"87",x"d1",x"e3"),
   495 => (x"31",x"c9",x"49",x"66"),
   496 => (x"66",x"c4",x"1e",x"71"),
   497 => (x"92",x"cc",x"c1",x"4a"),
   498 => (x"49",x"cc",x"ca",x"c3"),
   499 => (x"cb",x"fe",x"81",x"72"),
   500 => (x"f6",x"c2",x"87",x"fa"),
   501 => (x"66",x"c8",x"1e",x"e8"),
   502 => (x"92",x"cc",x"c1",x"4a"),
   503 => (x"49",x"cc",x"ca",x"c3"),
   504 => (x"c9",x"fe",x"81",x"72"),
   505 => (x"49",x"d7",x"87",x"e8"),
   506 => (x"87",x"f8",x"d8",x"ff"),
   507 => (x"c2",x"1e",x"c0",x"c8"),
   508 => (x"fd",x"49",x"e8",x"f6"),
   509 => (x"cc",x"87",x"d9",x"e4"),
   510 => (x"48",x"d0",x"ff",x"86"),
   511 => (x"f8",x"78",x"e0",x"c0"),
   512 => (x"26",x"4c",x"26",x"8e"),
   513 => (x"1e",x"4f",x"26",x"4b"),
   514 => (x"b7",x"c2",x"4a",x"71"),
   515 => (x"87",x"ce",x"03",x"aa"),
   516 => (x"cc",x"c1",x"49",x"72"),
   517 => (x"cc",x"ca",x"c3",x"91"),
   518 => (x"81",x"c8",x"c1",x"81"),
   519 => (x"4f",x"26",x"79",x"c0"),
   520 => (x"5c",x"5b",x"5e",x"0e"),
   521 => (x"86",x"fc",x"0e",x"5d"),
   522 => (x"d4",x"ff",x"4a",x"71"),
   523 => (x"d4",x"4c",x"c0",x"4b"),
   524 => (x"b7",x"c3",x"4d",x"66"),
   525 => (x"c2",x"c2",x"01",x"ad"),
   526 => (x"02",x"9a",x"72",x"87"),
   527 => (x"1e",x"87",x"ec",x"c0"),
   528 => (x"cc",x"c1",x"49",x"75"),
   529 => (x"cc",x"ca",x"c3",x"91"),
   530 => (x"c8",x"80",x"71",x"48"),
   531 => (x"66",x"c4",x"58",x"a6"),
   532 => (x"c3",x"c3",x"fe",x"49"),
   533 => (x"70",x"86",x"c4",x"87"),
   534 => (x"87",x"d4",x"02",x"98"),
   535 => (x"c8",x"c1",x"49",x"6e"),
   536 => (x"6e",x"79",x"c1",x"81"),
   537 => (x"69",x"81",x"c8",x"49"),
   538 => (x"75",x"87",x"c5",x"4c"),
   539 => (x"87",x"d7",x"fe",x"49"),
   540 => (x"c8",x"48",x"d0",x"ff"),
   541 => (x"7b",x"dd",x"78",x"e1"),
   542 => (x"ff",x"c3",x"48",x"74"),
   543 => (x"74",x"7b",x"70",x"98"),
   544 => (x"29",x"b7",x"c8",x"49"),
   545 => (x"ff",x"c3",x"48",x"71"),
   546 => (x"74",x"7b",x"70",x"98"),
   547 => (x"29",x"b7",x"d0",x"49"),
   548 => (x"ff",x"c3",x"48",x"71"),
   549 => (x"74",x"7b",x"70",x"98"),
   550 => (x"28",x"b7",x"d8",x"48"),
   551 => (x"7b",x"c0",x"7b",x"70"),
   552 => (x"7b",x"7b",x"7b",x"7b"),
   553 => (x"7b",x"7b",x"7b",x"7b"),
   554 => (x"ff",x"7b",x"7b",x"7b"),
   555 => (x"e0",x"c0",x"48",x"d0"),
   556 => (x"dc",x"1e",x"75",x"78"),
   557 => (x"d0",x"d6",x"ff",x"49"),
   558 => (x"fc",x"86",x"c4",x"87"),
   559 => (x"26",x"4d",x"26",x"8e"),
   560 => (x"26",x"4b",x"26",x"4c"),
   561 => (x"d4",x"ff",x"1e",x"4f"),
   562 => (x"7a",x"ff",x"c3",x"4a"),
   563 => (x"c5",x"48",x"d0",x"ff"),
   564 => (x"71",x"7a",x"c4",x"78"),
   565 => (x"28",x"b7",x"d8",x"48"),
   566 => (x"48",x"71",x"7a",x"70"),
   567 => (x"70",x"28",x"b7",x"d0"),
   568 => (x"c8",x"48",x"71",x"7a"),
   569 => (x"7a",x"70",x"28",x"b7"),
   570 => (x"d0",x"ff",x"7a",x"71"),
   571 => (x"26",x"78",x"c4",x"48"),
   572 => (x"4a",x"c0",x"1e",x"4f"),
   573 => (x"bf",x"e4",x"cc",x"c3"),
   574 => (x"49",x"87",x"ca",x"02"),
   575 => (x"48",x"e4",x"cc",x"c3"),
   576 => (x"11",x"78",x"a1",x"c1"),
   577 => (x"05",x"9a",x"72",x"4a"),
   578 => (x"cc",x"c3",x"87",x"c6"),
   579 => (x"78",x"c0",x"48",x"e4"),
   580 => (x"4f",x"26",x"48",x"72"),
   581 => (x"e4",x"cc",x"c3",x"1e"),
   582 => (x"c0",x"eb",x"c2",x"48"),
   583 => (x"4f",x"26",x"78",x"bf"),
   584 => (x"5c",x"5b",x"5e",x"0e"),
   585 => (x"ff",x"4a",x"71",x"0e"),
   586 => (x"d4",x"ff",x"4c",x"d0"),
   587 => (x"c1",x"7c",x"c5",x"4b"),
   588 => (x"7b",x"c3",x"7b",x"d5"),
   589 => (x"7c",x"c5",x"7c",x"c4"),
   590 => (x"c1",x"7b",x"d3",x"c1"),
   591 => (x"c8",x"7c",x"c4",x"7b"),
   592 => (x"d4",x"c1",x"7c",x"c5"),
   593 => (x"b7",x"49",x"c0",x"7b"),
   594 => (x"87",x"ca",x"06",x"aa"),
   595 => (x"81",x"c1",x"7b",x"c0"),
   596 => (x"04",x"a9",x"b7",x"72"),
   597 => (x"7c",x"c4",x"87",x"f6"),
   598 => (x"d3",x"c1",x"7c",x"c5"),
   599 => (x"c4",x"7b",x"c0",x"7b"),
   600 => (x"26",x"4c",x"26",x"7c"),
   601 => (x"1e",x"4f",x"26",x"4b"),
   602 => (x"4b",x"71",x"1e",x"73"),
   603 => (x"fc",x"c3",x"c3",x"1e"),
   604 => (x"e3",x"fe",x"fd",x"49"),
   605 => (x"70",x"86",x"c4",x"87"),
   606 => (x"e1",x"c0",x"02",x"98"),
   607 => (x"c4",x"c4",x"c3",x"87"),
   608 => (x"2a",x"ca",x"4a",x"bf"),
   609 => (x"02",x"8a",x"c0",x"c3"),
   610 => (x"c0",x"c1",x"87",x"ce"),
   611 => (x"87",x"ce",x"05",x"8a"),
   612 => (x"48",x"dc",x"e8",x"c1"),
   613 => (x"87",x"c6",x"50",x"c0"),
   614 => (x"48",x"dc",x"e8",x"c1"),
   615 => (x"4b",x"26",x"50",x"c1"),
   616 => (x"73",x"1e",x"4f",x"26"),
   617 => (x"f8",x"c3",x"c3",x"1e"),
   618 => (x"c1",x"50",x"c0",x"48"),
   619 => (x"c1",x"48",x"dc",x"e8"),
   620 => (x"c4",x"ff",x"c0",x"50"),
   621 => (x"c1",x"50",x"c0",x"48"),
   622 => (x"87",x"c9",x"fc",x"49"),
   623 => (x"49",x"c0",x"c0",x"c4"),
   624 => (x"c2",x"87",x"dd",x"fd"),
   625 => (x"49",x"bf",x"d4",x"eb"),
   626 => (x"c2",x"87",x"dc",x"fe"),
   627 => (x"49",x"bf",x"d4",x"eb"),
   628 => (x"87",x"d6",x"d8",x"fe"),
   629 => (x"ec",x"fb",x"49",x"c0"),
   630 => (x"49",x"d0",x"c6",x"87"),
   631 => (x"70",x"87",x"f1",x"f2"),
   632 => (x"f7",x"f2",x"49",x"4b"),
   633 => (x"05",x"98",x"70",x"87"),
   634 => (x"49",x"73",x"87",x"ca"),
   635 => (x"70",x"87",x"ed",x"f2"),
   636 => (x"87",x"f6",x"02",x"98"),
   637 => (x"cc",x"fb",x"49",x"c1"),
   638 => (x"49",x"e4",x"c1",x"87"),
   639 => (x"70",x"87",x"d1",x"f2"),
   640 => (x"d7",x"f2",x"49",x"4b"),
   641 => (x"05",x"98",x"70",x"87"),
   642 => (x"49",x"73",x"87",x"ca"),
   643 => (x"70",x"87",x"cd",x"f2"),
   644 => (x"87",x"f6",x"02",x"98"),
   645 => (x"ec",x"fa",x"49",x"c0"),
   646 => (x"26",x"48",x"c0",x"87"),
   647 => (x"1e",x"4f",x"26",x"4b"),
   648 => (x"ea",x"c2",x"1e",x"73"),
   649 => (x"c0",x"05",x"bf",x"fc"),
   650 => (x"c9",x"c3",x"87",x"ea"),
   651 => (x"c4",x"ff",x"49",x"d8"),
   652 => (x"b7",x"c0",x"87",x"e8"),
   653 => (x"87",x"ce",x"04",x"a8"),
   654 => (x"49",x"d8",x"c9",x"c3"),
   655 => (x"87",x"da",x"c4",x"ff"),
   656 => (x"03",x"a8",x"b7",x"c0"),
   657 => (x"ea",x"c2",x"87",x"f2"),
   658 => (x"c1",x"48",x"bf",x"fc"),
   659 => (x"c0",x"eb",x"c2",x"80"),
   660 => (x"87",x"e2",x"c1",x"58"),
   661 => (x"bf",x"fc",x"ea",x"c2"),
   662 => (x"99",x"c1",x"49",x"4b"),
   663 => (x"87",x"f0",x"c0",x"02"),
   664 => (x"b7",x"c1",x"49",x"73"),
   665 => (x"d8",x"eb",x"c2",x"29"),
   666 => (x"9a",x"4a",x"11",x"81"),
   667 => (x"87",x"c6",x"c1",x"02"),
   668 => (x"06",x"aa",x"b7",x"c1"),
   669 => (x"1e",x"72",x"87",x"cc"),
   670 => (x"49",x"d8",x"c9",x"c3"),
   671 => (x"87",x"e6",x"c1",x"ff"),
   672 => (x"ea",x"c2",x"86",x"c4"),
   673 => (x"c1",x"48",x"bf",x"fc"),
   674 => (x"c0",x"eb",x"c2",x"80"),
   675 => (x"87",x"e6",x"c0",x"58"),
   676 => (x"49",x"d8",x"c9",x"c3"),
   677 => (x"87",x"c2",x"c3",x"ff"),
   678 => (x"ea",x"c2",x"4a",x"70"),
   679 => (x"87",x"cb",x"02",x"aa"),
   680 => (x"02",x"aa",x"fa",x"c3"),
   681 => (x"aa",x"c3",x"87",x"c5"),
   682 => (x"c2",x"87",x"cb",x"05"),
   683 => (x"48",x"bf",x"fc",x"ea"),
   684 => (x"eb",x"c2",x"80",x"c1"),
   685 => (x"4b",x"26",x"58",x"c0"),
   686 => (x"00",x"00",x"4f",x"26"),
   687 => (x"00",x"00",x"00",x"00"),
   688 => (x"00",x"00",x"2b",x"f0"),
   689 => (x"11",x"14",x"12",x"58"),
   690 => (x"23",x"1c",x"1b",x"1d"),
   691 => (x"91",x"94",x"59",x"5a"),
   692 => (x"f4",x"eb",x"f2",x"f5"),
   693 => (x"00",x"00",x"2d",x"68"),
   694 => (x"f3",x"c8",x"f3",x"ff"),
   695 => (x"f2",x"50",x"f3",x"64"),
   696 => (x"1e",x"00",x"f4",x"01"),
   697 => (x"4b",x"71",x"1e",x"73"),
   698 => (x"c5",x"e8",x"fe",x"49"),
   699 => (x"fc",x"c9",x"c3",x"87"),
   700 => (x"c7",x"02",x"bf",x"97"),
   701 => (x"c0",x"c0",x"c4",x"87"),
   702 => (x"87",x"e4",x"f8",x"49"),
   703 => (x"e7",x"fe",x"49",x"73"),
   704 => (x"4b",x"26",x"87",x"f0"),
   705 => (x"73",x"1e",x"4f",x"26"),
   706 => (x"c3",x"4a",x"71",x"1e"),
   707 => (x"4b",x"bf",x"f0",x"c3"),
   708 => (x"c5",x"02",x"9a",x"72"),
   709 => (x"bb",x"c0",x"c2",x"87"),
   710 => (x"c0",x"c1",x"87",x"c3"),
   711 => (x"f6",x"49",x"73",x"bb"),
   712 => (x"f4",x"c7",x"87",x"e3"),
   713 => (x"87",x"e8",x"ed",x"49"),
   714 => (x"ed",x"49",x"4b",x"70"),
   715 => (x"98",x"70",x"87",x"ee"),
   716 => (x"73",x"87",x"ca",x"05"),
   717 => (x"87",x"e4",x"ed",x"49"),
   718 => (x"f6",x"02",x"98",x"70"),
   719 => (x"26",x"4b",x"26",x"87"),
   720 => (x"5b",x"5e",x"0e",x"4f"),
   721 => (x"4b",x"71",x"0e",x"5c"),
   722 => (x"d3",x"02",x"66",x"cc"),
   723 => (x"f0",x"c0",x"4c",x"87"),
   724 => (x"e9",x"c0",x"02",x"8c"),
   725 => (x"c1",x"49",x"74",x"87"),
   726 => (x"e1",x"c0",x"02",x"89"),
   727 => (x"87",x"f3",x"c0",x"87"),
   728 => (x"c0",x"02",x"9b",x"73"),
   729 => (x"c3",x"c3",x"87",x"ed"),
   730 => (x"c1",x"49",x"bf",x"f0"),
   731 => (x"d4",x"f5",x"71",x"b1"),
   732 => (x"f7",x"49",x"73",x"87"),
   733 => (x"49",x"73",x"87",x"f1"),
   734 => (x"87",x"ee",x"d1",x"fe"),
   735 => (x"1e",x"74",x"87",x"d5"),
   736 => (x"db",x"f2",x"49",x"c0"),
   737 => (x"fd",x"49",x"74",x"87"),
   738 => (x"1e",x"74",x"87",x"fc"),
   739 => (x"cf",x"f2",x"49",x"73"),
   740 => (x"c3",x"86",x"c8",x"87"),
   741 => (x"49",x"bf",x"f0",x"c3"),
   742 => (x"26",x"87",x"ea",x"f4"),
   743 => (x"26",x"4b",x"26",x"4c"),
   744 => (x"c4",x"ff",x"1e",x"4f"),
   745 => (x"d4",x"ff",x"87",x"df"),
   746 => (x"78",x"ff",x"c3",x"48"),
   747 => (x"87",x"d0",x"df",x"fd"),
   748 => (x"cd",x"02",x"98",x"70"),
   749 => (x"ee",x"e8",x"fd",x"87"),
   750 => (x"02",x"98",x"70",x"87"),
   751 => (x"4a",x"c1",x"87",x"c4"),
   752 => (x"4a",x"c0",x"87",x"c2"),
   753 => (x"c8",x"02",x"9a",x"72"),
   754 => (x"ec",x"ef",x"c2",x"87"),
   755 => (x"d6",x"d3",x"fd",x"49"),
   756 => (x"fe",x"49",x"c0",x"87"),
   757 => (x"f7",x"87",x"e1",x"f8"),
   758 => (x"fb",x"fe",x"87",x"c8"),
   759 => (x"fe",x"f8",x"87",x"e1"),
   760 => (x"e5",x"de",x"ff",x"87"),
   761 => (x"87",x"c1",x"ed",x"87"),
   762 => (x"4f",x"26",x"87",x"f4"),
   763 => (x"00",x"00",x"4b",x"4f"),
   764 => (x"72",x"61",x"74",x"41"),
   765 => (x"54",x"53",x"20",x"69"),
   766 => (x"30",x"53",x"3b",x"3b"),
   767 => (x"54",x"53",x"2c",x"55"),
   768 => (x"6c",x"46",x"2c",x"20"),
   769 => (x"79",x"70",x"70",x"6f"),
   770 => (x"3b",x"3a",x"41",x"20"),
   771 => (x"2c",x"55",x"31",x"53"),
   772 => (x"2c",x"20",x"54",x"53"),
   773 => (x"70",x"6f",x"6c",x"46"),
   774 => (x"42",x"20",x"79",x"70"),
   775 => (x"36",x"4f",x"3b",x"3a"),
   776 => (x"72",x"57",x"2c",x"37"),
   777 => (x"20",x"65",x"74",x"69"),
   778 => (x"74",x"6f",x"72",x"70"),
   779 => (x"2c",x"74",x"63",x"65"),
   780 => (x"2c",x"66",x"66",x"4f"),
   781 => (x"42",x"2c",x"3a",x"41"),
   782 => (x"6f",x"42",x"2c",x"3a"),
   783 => (x"46",x"3b",x"68",x"74"),
   784 => (x"47",x"4d",x"49",x"2c"),
   785 => (x"2c",x"4d",x"4f",x"52"),
   786 => (x"64",x"61",x"6f",x"4c"),
   787 => (x"4d",x"4f",x"52",x"20"),
   788 => (x"2c",x"31",x"50",x"3b"),
   789 => (x"43",x"20",x"54",x"53"),
   790 => (x"69",x"66",x"6e",x"6f"),
   791 => (x"61",x"72",x"75",x"67"),
   792 => (x"6e",x"6f",x"69",x"74"),
   793 => (x"4f",x"31",x"50",x"3b"),
   794 => (x"52",x"2c",x"33",x"31"),
   795 => (x"28",x"20",x"4d",x"41"),
   796 => (x"64",x"65",x"65",x"6e"),
   797 => (x"72",x"61",x"48",x"20"),
   798 => (x"65",x"52",x"20",x"64"),
   799 => (x"29",x"74",x"65",x"73"),
   800 => (x"32",x"31",x"35",x"2c"),
   801 => (x"4d",x"31",x"2c",x"4b"),
   802 => (x"4d",x"32",x"2c",x"42"),
   803 => (x"4d",x"34",x"2c",x"42"),
   804 => (x"4d",x"38",x"2c",x"42"),
   805 => (x"34",x"31",x"2c",x"42"),
   806 => (x"50",x"3b",x"42",x"4d"),
   807 => (x"2c",x"38",x"4f",x"31"),
   808 => (x"65",x"64",x"69",x"56"),
   809 => (x"6f",x"6d",x"20",x"6f"),
   810 => (x"4d",x"2c",x"65",x"64"),
   811 => (x"2c",x"6f",x"6e",x"6f"),
   812 => (x"6f",x"6c",x"6f",x"43"),
   813 => (x"50",x"3b",x"72",x"75"),
   814 => (x"4f",x"4e",x"4f",x"31"),
   815 => (x"69",x"68",x"43",x"2c"),
   816 => (x"74",x"65",x"73",x"70"),
   817 => (x"2c",x"54",x"53",x"2c"),
   818 => (x"2c",x"45",x"54",x"53"),
   819 => (x"61",x"67",x"65",x"4d"),
   820 => (x"3b",x"45",x"54",x"53"),
   821 => (x"4a",x"4f",x"31",x"50"),
   822 => (x"20",x"54",x"53",x"2c"),
   823 => (x"74",x"69",x"6c",x"42"),
   824 => (x"2c",x"72",x"65",x"74"),
   825 => (x"2c",x"66",x"66",x"4f"),
   826 => (x"50",x"3b",x"6e",x"4f"),
   827 => (x"2c",x"4d",x"4f",x"31"),
   828 => (x"72",x"65",x"74",x"53"),
   829 => (x"73",x"20",x"6f",x"65"),
   830 => (x"64",x"6e",x"75",x"6f"),
   831 => (x"66",x"66",x"4f",x"2c"),
   832 => (x"3b",x"6e",x"4f",x"2c"),
   833 => (x"4b",x"4f",x"31",x"50"),
   834 => (x"63",x"53",x"2c",x"4c"),
   835 => (x"69",x"6c",x"6e",x"61"),
   836 => (x"2c",x"73",x"65",x"6e"),
   837 => (x"2c",x"66",x"66",x"4f"),
   838 => (x"2c",x"25",x"35",x"32"),
   839 => (x"2c",x"25",x"30",x"35"),
   840 => (x"3b",x"25",x"35",x"37"),
   841 => (x"54",x"4f",x"31",x"50"),
   842 => (x"6d",x"6f",x"43",x"2c"),
   843 => (x"69",x"73",x"6f",x"70"),
   844 => (x"62",x"20",x"65",x"74"),
   845 => (x"64",x"6e",x"65",x"6c"),
   846 => (x"66",x"66",x"4f",x"2c"),
   847 => (x"3b",x"6e",x"4f",x"2c"),
   848 => (x"52",x"2c",x"30",x"54"),
   849 => (x"74",x"65",x"73",x"65"),
   850 => (x"6f",x"48",x"28",x"20"),
   851 => (x"66",x"20",x"64",x"6c"),
   852 => (x"68",x"20",x"72",x"6f"),
   853 => (x"20",x"64",x"72",x"61"),
   854 => (x"65",x"73",x"65",x"72"),
   855 => (x"56",x"3b",x"29",x"74"),
   856 => (x"2e",x"33",x"76",x"2c"),
   857 => (x"00",x"2e",x"30",x"34"),
   858 => (x"20",x"53",x"4f",x"54"),
   859 => (x"20",x"20",x"20",x"20"),
   860 => (x"00",x"47",x"4d",x"49"),
   861 => (x"00",x"00",x"1a",x"af"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

