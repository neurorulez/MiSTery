library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e8ccc387",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49e8ccc3",
    18 => x"48f8f5c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"f8f5c287",
    25 => x"f4f5c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"ecc287f7",
    29 => x"f5c287eb",
    30 => x"f5c24df8",
    31 => x"ad744cf8",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"8148731e",
    65 => x"c502a973",
    66 => x"05531287",
    67 => x"4f2687f6",
    68 => x"711e731e",
    69 => x"4b66c84a",
    70 => x"718bc149",
    71 => x"87cf0299",
    72 => x"d4ff4812",
    73 => x"49737808",
    74 => x"99718bc1",
    75 => x"2687f105",
    76 => x"0e4f264b",
    77 => x"0e5c5b5e",
    78 => x"d4ff4a71",
    79 => x"4b66cc4c",
    80 => x"718bc149",
    81 => x"87ce0299",
    82 => x"6c7cffc3",
    83 => x"c1497352",
    84 => x"0599718b",
    85 => x"4c2687f2",
    86 => x"4f264b26",
    87 => x"ff1e731e",
    88 => x"ffc34bd4",
    89 => x"c34a6b7b",
    90 => x"496b7bff",
    91 => x"b17232c8",
    92 => x"6b7bffc3",
    93 => x"7131c84a",
    94 => x"7bffc3b2",
    95 => x"32c8496b",
    96 => x"4871b172",
    97 => x"4f264b26",
    98 => x"5c5b5e0e",
    99 => x"4d710e5d",
   100 => x"754cd4ff",
   101 => x"98ffc348",
   102 => x"f5c27c70",
   103 => x"c805bff8",
   104 => x"4866d087",
   105 => x"a6d430c9",
   106 => x"4966d058",
   107 => x"487129d8",
   108 => x"7098ffc3",
   109 => x"4966d07c",
   110 => x"487129d0",
   111 => x"7098ffc3",
   112 => x"4966d07c",
   113 => x"487129c8",
   114 => x"7098ffc3",
   115 => x"4866d07c",
   116 => x"7098ffc3",
   117 => x"d049757c",
   118 => x"c3487129",
   119 => x"7c7098ff",
   120 => x"f0c94b6c",
   121 => x"ffc34aff",
   122 => x"87cf05ab",
   123 => x"6c7c7149",
   124 => x"028ac14b",
   125 => x"ab7187c5",
   126 => x"7387f202",
   127 => x"264d2648",
   128 => x"264b264c",
   129 => x"49c01e4f",
   130 => x"c348d4ff",
   131 => x"81c178ff",
   132 => x"a9b7c8c3",
   133 => x"2687f104",
   134 => x"5b5e0e4f",
   135 => x"c00e5d5c",
   136 => x"f7c1f0ff",
   137 => x"c0c0c14d",
   138 => x"4bc0c0c0",
   139 => x"c487d6ff",
   140 => x"c04cdff8",
   141 => x"fd49751e",
   142 => x"86c487ce",
   143 => x"c005a8c1",
   144 => x"d4ff87e5",
   145 => x"78ffc348",
   146 => x"e1c01e73",
   147 => x"49e9c1f0",
   148 => x"c487f5fc",
   149 => x"05987086",
   150 => x"d4ff87ca",
   151 => x"78ffc348",
   152 => x"87cb48c1",
   153 => x"c187defe",
   154 => x"c6ff058c",
   155 => x"2648c087",
   156 => x"264c264d",
   157 => x"0e4f264b",
   158 => x"0e5c5b5e",
   159 => x"c1f0ffc0",
   160 => x"d4ff4cc1",
   161 => x"78ffc348",
   162 => x"f849fcca",
   163 => x"4bd387d9",
   164 => x"49741ec0",
   165 => x"c487f1fb",
   166 => x"05987086",
   167 => x"d4ff87ca",
   168 => x"78ffc348",
   169 => x"87cb48c1",
   170 => x"c187dafd",
   171 => x"dfff058b",
   172 => x"2648c087",
   173 => x"264b264c",
   174 => x"0000004f",
   175 => x"00444d43",
   176 => x"43484453",
   177 => x"69616620",
   178 => x"000a216c",
   179 => x"52524549",
   180 => x"00000000",
   181 => x"00495053",
   182 => x"74697257",
   183 => x"61662065",
   184 => x"64656c69",
   185 => x"5e0e000a",
   186 => x"0e5d5c5b",
   187 => x"ff4dffc3",
   188 => x"d0fc4bd4",
   189 => x"1eeac687",
   190 => x"c1f0e1c0",
   191 => x"c7fa49c8",
   192 => x"c186c487",
   193 => x"87c802a8",
   194 => x"c087ecfd",
   195 => x"87e8c148",
   196 => x"7087c9f9",
   197 => x"ffffcf49",
   198 => x"a9eac699",
   199 => x"fd87c802",
   200 => x"48c087d5",
   201 => x"7587d1c1",
   202 => x"4cf1c07b",
   203 => x"7087eafb",
   204 => x"ecc00298",
   205 => x"c01ec087",
   206 => x"fac1f0ff",
   207 => x"87c8f949",
   208 => x"987086c4",
   209 => x"7587da05",
   210 => x"75496b7b",
   211 => x"757b757b",
   212 => x"c17b757b",
   213 => x"c40299c0",
   214 => x"db48c187",
   215 => x"d748c087",
   216 => x"05acc287",
   217 => x"c0cb87ca",
   218 => x"87fbf449",
   219 => x"87c848c0",
   220 => x"fe058cc1",
   221 => x"48c087f6",
   222 => x"4c264d26",
   223 => x"4f264b26",
   224 => x"5c5b5e0e",
   225 => x"d0ff0e5d",
   226 => x"d0e5c04d",
   227 => x"c24cc0c1",
   228 => x"c148f8f5",
   229 => x"49d4cb78",
   230 => x"c787ccf4",
   231 => x"f97dc24b",
   232 => x"7dc387e3",
   233 => x"49741ec0",
   234 => x"c487ddf7",
   235 => x"05a8c186",
   236 => x"c24b87c1",
   237 => x"87cb05ab",
   238 => x"f349cccb",
   239 => x"48c087e9",
   240 => x"c187f6c0",
   241 => x"d4ff058b",
   242 => x"87dafc87",
   243 => x"58fcf5c2",
   244 => x"cd059870",
   245 => x"c01ec187",
   246 => x"d0c1f0ff",
   247 => x"87e8f649",
   248 => x"d4ff86c4",
   249 => x"78ffc348",
   250 => x"c287eec4",
   251 => x"c258c0f6",
   252 => x"48d4ff7d",
   253 => x"c178ffc3",
   254 => x"264d2648",
   255 => x"264b264c",
   256 => x"5b5e0e4f",
   257 => x"710e5d5c",
   258 => x"4cffc34d",
   259 => x"744bd4ff",
   260 => x"48d0ff7b",
   261 => x"7478c3c4",
   262 => x"c01e757b",
   263 => x"d8c1f0ff",
   264 => x"87e4f549",
   265 => x"987086c4",
   266 => x"cb87cb02",
   267 => x"f6f149d8",
   268 => x"c048c187",
   269 => x"7b7487ee",
   270 => x"c87bfec3",
   271 => x"66d41ec0",
   272 => x"87ccf349",
   273 => x"7b7486c4",
   274 => x"7b747b74",
   275 => x"4ae0dad8",
   276 => x"056b7b74",
   277 => x"8ac187c5",
   278 => x"7487f505",
   279 => x"48d0ff7b",
   280 => x"48c078c2",
   281 => x"4c264d26",
   282 => x"4f264b26",
   283 => x"5c5b5e0e",
   284 => x"86fc0e5d",
   285 => x"d4ff4b71",
   286 => x"c57ec04c",
   287 => x"4adfcdee",
   288 => x"6c7cffc3",
   289 => x"a8fec348",
   290 => x"87f8c005",
   291 => x"9b734d74",
   292 => x"d487cc02",
   293 => x"49731e66",
   294 => x"c487d8f2",
   295 => x"ff87d486",
   296 => x"d1c448d0",
   297 => x"4a66d478",
   298 => x"c17dffc3",
   299 => x"87f8058a",
   300 => x"c35aa6d8",
   301 => x"737c7cff",
   302 => x"87c5059b",
   303 => x"d048d0ff",
   304 => x"7e4ac178",
   305 => x"fe058ac1",
   306 => x"486e87f6",
   307 => x"4d268efc",
   308 => x"4b264c26",
   309 => x"731e4f26",
   310 => x"c04a711e",
   311 => x"48d4ff4b",
   312 => x"ff78ffc3",
   313 => x"c3c448d0",
   314 => x"48d4ff78",
   315 => x"7278ffc3",
   316 => x"f0ffc01e",
   317 => x"f249d1c1",
   318 => x"86c487ce",
   319 => x"d2059870",
   320 => x"1ec0c887",
   321 => x"fd4966cc",
   322 => x"86c487e2",
   323 => x"d0ff4b70",
   324 => x"7378c248",
   325 => x"264b2648",
   326 => x"5b5e0e4f",
   327 => x"c00e5d5c",
   328 => x"f0ffc01e",
   329 => x"f149c9c1",
   330 => x"1ed287de",
   331 => x"49c8f6c2",
   332 => x"c887f9fc",
   333 => x"c14cc086",
   334 => x"acb7d284",
   335 => x"c287f804",
   336 => x"bf97c8f6",
   337 => x"99c0c349",
   338 => x"05a9c0c1",
   339 => x"c287e7c0",
   340 => x"bf97cff6",
   341 => x"c231d049",
   342 => x"bf97d0f6",
   343 => x"7232c84a",
   344 => x"d1f6c2b1",
   345 => x"b14abf97",
   346 => x"ffcf4c71",
   347 => x"c19cffff",
   348 => x"c134ca84",
   349 => x"f6c287e7",
   350 => x"49bf97d1",
   351 => x"99c631c1",
   352 => x"97d2f6c2",
   353 => x"b7c74abf",
   354 => x"c2b1722a",
   355 => x"bf97cdf6",
   356 => x"9dcf4d4a",
   357 => x"97cef6c2",
   358 => x"9ac34abf",
   359 => x"f6c232ca",
   360 => x"4bbf97cf",
   361 => x"b27333c2",
   362 => x"97d0f6c2",
   363 => x"c0c34bbf",
   364 => x"2bb7c69b",
   365 => x"81c2b273",
   366 => x"307148c1",
   367 => x"48c14970",
   368 => x"4d703075",
   369 => x"84c14c72",
   370 => x"c0c89471",
   371 => x"cc06adb7",
   372 => x"b734c187",
   373 => x"b7c0c82d",
   374 => x"f4ff01ad",
   375 => x"26487487",
   376 => x"264c264d",
   377 => x"0e4f264b",
   378 => x"5d5c5b5e",
   379 => x"c286fc0e",
   380 => x"c048f0fe",
   381 => x"e8f6c278",
   382 => x"fb49c01e",
   383 => x"86c487d8",
   384 => x"c5059870",
   385 => x"c948c087",
   386 => x"4dc087d2",
   387 => x"48ecc3c3",
   388 => x"f7c278c1",
   389 => x"e1c04ade",
   390 => x"4bc849f4",
   391 => x"7087c7eb",
   392 => x"87c60598",
   393 => x"48ecc3c3",
   394 => x"f7c278c0",
   395 => x"e2c04afa",
   396 => x"4bc849c0",
   397 => x"7087efea",
   398 => x"87c60598",
   399 => x"48ecc3c3",
   400 => x"c3c378c0",
   401 => x"c002bfec",
   402 => x"fdc287fd",
   403 => x"c24dbfee",
   404 => x"bf9fe6fe",
   405 => x"d6c5487e",
   406 => x"c705a8ea",
   407 => x"eefdc287",
   408 => x"87ce4dbf",
   409 => x"e9ca486e",
   410 => x"c502a8d5",
   411 => x"c748c087",
   412 => x"f6c287ea",
   413 => x"49751ee8",
   414 => x"c487dbf9",
   415 => x"05987086",
   416 => x"48c087c5",
   417 => x"c287d5c7",
   418 => x"c04afaf7",
   419 => x"c849cce2",
   420 => x"87d2e94b",
   421 => x"c8059870",
   422 => x"f0fec287",
   423 => x"d878c148",
   424 => x"def7c287",
   425 => x"d8e2c04a",
   426 => x"e84bc849",
   427 => x"987087f8",
   428 => x"87c5c002",
   429 => x"e3c648c0",
   430 => x"e6fec287",
   431 => x"c149bf97",
   432 => x"c005a9d5",
   433 => x"fec287cd",
   434 => x"49bf97e7",
   435 => x"02a9eac2",
   436 => x"c087c5c0",
   437 => x"87c4c648",
   438 => x"97e8f6c2",
   439 => x"c3487ebf",
   440 => x"c002a8e9",
   441 => x"486e87ce",
   442 => x"02a8ebc3",
   443 => x"c087c5c0",
   444 => x"87e8c548",
   445 => x"97f3f6c2",
   446 => x"059949bf",
   447 => x"c287ccc0",
   448 => x"bf97f4f6",
   449 => x"02a9c249",
   450 => x"c087c5c0",
   451 => x"87ccc548",
   452 => x"97f5f6c2",
   453 => x"fec248bf",
   454 => x"4c7058ec",
   455 => x"c288c148",
   456 => x"c258f0fe",
   457 => x"bf97f6f6",
   458 => x"c2817549",
   459 => x"bf97f7f6",
   460 => x"7232c84a",
   461 => x"c3c37ea1",
   462 => x"786e48c8",
   463 => x"97f8f6c2",
   464 => x"c3c348bf",
   465 => x"fec258e0",
   466 => x"c202bff0",
   467 => x"f7c287d3",
   468 => x"e1c04afa",
   469 => x"4bc849e8",
   470 => x"7087cbe6",
   471 => x"c5c00298",
   472 => x"c348c087",
   473 => x"fec287f6",
   474 => x"c34cbfe8",
   475 => x"c25cdcc3",
   476 => x"bf97cdf7",
   477 => x"c231c849",
   478 => x"bf97ccf7",
   479 => x"c249a14a",
   480 => x"bf97cef7",
   481 => x"7232d04a",
   482 => x"f7c249a1",
   483 => x"4abf97cf",
   484 => x"a17232d8",
   485 => x"e4c3c349",
   486 => x"dcc3c359",
   487 => x"c3c391bf",
   488 => x"c381bfc8",
   489 => x"c259d0c3",
   490 => x"bf97d5f7",
   491 => x"c232c84a",
   492 => x"bf97d4f7",
   493 => x"c24aa24b",
   494 => x"bf97d6f7",
   495 => x"7333d04b",
   496 => x"f7c24aa2",
   497 => x"4bbf97d7",
   498 => x"33d89bcf",
   499 => x"c34aa273",
   500 => x"c25ad4c3",
   501 => x"c392748a",
   502 => x"7248d4c3",
   503 => x"c7c178a1",
   504 => x"faf6c287",
   505 => x"c849bf97",
   506 => x"f9f6c231",
   507 => x"a14abf97",
   508 => x"c731c549",
   509 => x"29c981ff",
   510 => x"59dcc3c3",
   511 => x"97fff6c2",
   512 => x"32c84abf",
   513 => x"97fef6c2",
   514 => x"4aa24bbf",
   515 => x"5ae4c3c3",
   516 => x"bfdcc3c3",
   517 => x"c3826e92",
   518 => x"c35ad8c3",
   519 => x"c048d0c3",
   520 => x"ccc3c378",
   521 => x"78a17248",
   522 => x"48e4c3c3",
   523 => x"bfd0c3c3",
   524 => x"e8c3c378",
   525 => x"d4c3c348",
   526 => x"fec278bf",
   527 => x"c002bff0",
   528 => x"487487c9",
   529 => x"7e7030c4",
   530 => x"c387c9c0",
   531 => x"48bfd8c3",
   532 => x"7e7030c4",
   533 => x"48f4fec2",
   534 => x"48c1786e",
   535 => x"4d268efc",
   536 => x"4b264c26",
   537 => x"00004f26",
   538 => x"33544146",
   539 => x"20202032",
   540 => x"00000000",
   541 => x"31544146",
   542 => x"20202036",
   543 => x"00000000",
   544 => x"33544146",
   545 => x"20202032",
   546 => x"00000000",
   547 => x"33544146",
   548 => x"20202032",
   549 => x"00000000",
   550 => x"31544146",
   551 => x"20202036",
   552 => x"5b5e0e00",
   553 => x"710e5d5c",
   554 => x"f0fec24a",
   555 => x"87cb02bf",
   556 => x"2bc74b72",
   557 => x"ffc14d72",
   558 => x"7287c99d",
   559 => x"722bc84b",
   560 => x"9dffc34d",
   561 => x"bfc8c3c3",
   562 => x"e8f9c083",
   563 => x"d902abbf",
   564 => x"ecf9c087",
   565 => x"e8f6c25b",
   566 => x"ef49731e",
   567 => x"86c487f8",
   568 => x"c5059870",
   569 => x"c048c087",
   570 => x"fec287e6",
   571 => x"d202bff0",
   572 => x"c4497587",
   573 => x"e8f6c291",
   574 => x"cf4c6981",
   575 => x"ffffffff",
   576 => x"7587cb9c",
   577 => x"c291c249",
   578 => x"9f81e8f6",
   579 => x"48744c69",
   580 => x"4c264d26",
   581 => x"4f264b26",
   582 => x"5c5b5e0e",
   583 => x"86f40e5d",
   584 => x"c459a6c8",
   585 => x"80c84866",
   586 => x"c0487e70",
   587 => x"49c11e78",
   588 => x"87f9cc49",
   589 => x"4c7086c4",
   590 => x"fcc0029c",
   591 => x"f8fec287",
   592 => x"4966dc4a",
   593 => x"87c3deff",
   594 => x"c0029870",
   595 => x"4a7487eb",
   596 => x"cb4966dc",
   597 => x"cddeff4b",
   598 => x"02987087",
   599 => x"1ec087db",
   600 => x"c4029c74",
   601 => x"c24dc087",
   602 => x"754dc187",
   603 => x"87fdcb49",
   604 => x"4c7086c4",
   605 => x"c4ff059c",
   606 => x"029c7487",
   607 => x"dc87f4c1",
   608 => x"486e49a4",
   609 => x"a4da7869",
   610 => x"4d66c449",
   611 => x"699f85c4",
   612 => x"f0fec27d",
   613 => x"87d202bf",
   614 => x"9f49a4d4",
   615 => x"ffc04969",
   616 => x"487199ff",
   617 => x"7e7030d0",
   618 => x"7ec087c2",
   619 => x"6d48496e",
   620 => x"c47d7080",
   621 => x"78c04866",
   622 => x"cc4966c4",
   623 => x"c4796d81",
   624 => x"81d04966",
   625 => x"a6c879c0",
   626 => x"c878c048",
   627 => x"66c44c66",
   628 => x"7482d44a",
   629 => x"7291c849",
   630 => x"41c049a1",
   631 => x"84c1796d",
   632 => x"04acb7c6",
   633 => x"c487e7ff",
   634 => x"c4c14966",
   635 => x"c179c081",
   636 => x"c087c248",
   637 => x"268ef448",
   638 => x"264c264d",
   639 => x"0e4f264b",
   640 => x"5d5c5b5e",
   641 => x"d04c710e",
   642 => x"6c4a4d66",
   643 => x"4da17249",
   644 => x"ecfec2b9",
   645 => x"baff4abf",
   646 => x"99719972",
   647 => x"87e4c002",
   648 => x"6b4ba4c4",
   649 => x"87f9f949",
   650 => x"fec27b70",
   651 => x"6c49bfe8",
   652 => x"757c7181",
   653 => x"ecfec2b9",
   654 => x"baff4abf",
   655 => x"99719972",
   656 => x"87dcff05",
   657 => x"4d267c75",
   658 => x"4b264c26",
   659 => x"731e4f26",
   660 => x"c34b711e",
   661 => x"49bfccc3",
   662 => x"6a4aa3c4",
   663 => x"c28ac24a",
   664 => x"92bfe8fe",
   665 => x"c249a172",
   666 => x"4abfecfe",
   667 => x"a1729a6b",
   668 => x"ecf9c049",
   669 => x"1e66c859",
   670 => x"87dae971",
   671 => x"987086c4",
   672 => x"c087c405",
   673 => x"c187c248",
   674 => x"264b2648",
   675 => x"1e731e4f",
   676 => x"c3c34b71",
   677 => x"c449bfcc",
   678 => x"4a6a4aa3",
   679 => x"fec28ac2",
   680 => x"7292bfe8",
   681 => x"fec249a1",
   682 => x"6b4abfec",
   683 => x"49a1729a",
   684 => x"59ecf9c0",
   685 => x"711e66c8",
   686 => x"c487c6e5",
   687 => x"05987086",
   688 => x"48c087c4",
   689 => x"48c187c2",
   690 => x"4f264b26",
   691 => x"5c5b5e0e",
   692 => x"86e00e5d",
   693 => x"f0c04b71",
   694 => x"29c94966",
   695 => x"c259a6c8",
   696 => x"49bfecfe",
   697 => x"4a71b9ff",
   698 => x"d89a66c4",
   699 => x"996b5aa6",
   700 => x"c459a6d0",
   701 => x"a6d07ea3",
   702 => x"78bf6e48",
   703 => x"cc4866d4",
   704 => x"c605a866",
   705 => x"7b66c487",
   706 => x"d887c1c3",
   707 => x"ffc148a6",
   708 => x"ffffffff",
   709 => x"ff80c478",
   710 => x"c84cc078",
   711 => x"a3d448a6",
   712 => x"c8497478",
   713 => x"8166c891",
   714 => x"4d4a66d4",
   715 => x"b7c08d69",
   716 => x"87ce04ad",
   717 => x"adb766d8",
   718 => x"c087c703",
   719 => x"dc5ca6e0",
   720 => x"84c15da6",
   721 => x"04acb7c6",
   722 => x"dc87d0ff",
   723 => x"b7c04866",
   724 => x"87d004a8",
   725 => x"c84966dc",
   726 => x"8166c891",
   727 => x"486e7b21",
   728 => x"87c97869",
   729 => x"a3cc7bc0",
   730 => x"69486e49",
   731 => x"4866c478",
   732 => x"a6c8886b",
   733 => x"e8fec258",
   734 => x"90c848bf",
   735 => x"66c47e70",
   736 => x"01a86e48",
   737 => x"66c487c9",
   738 => x"03a86e48",
   739 => x"c187f3c0",
   740 => x"6a4aa3c4",
   741 => x"c891c849",
   742 => x"66cc8166",
   743 => x"c8496a79",
   744 => x"8166c891",
   745 => x"66d081c4",
   746 => x"487e6a79",
   747 => x"c705a8c5",
   748 => x"48a6c887",
   749 => x"87c778c0",
   750 => x"80c1486e",
   751 => x"c858a6cc",
   752 => x"66c47a66",
   753 => x"f849731e",
   754 => x"86c487f5",
   755 => x"1ee8f6c2",
   756 => x"f9f94973",
   757 => x"49a3d087",
   758 => x"7966f4c0",
   759 => x"268edcff",
   760 => x"264c264d",
   761 => x"0e4f264b",
   762 => x"0e5c5b5e",
   763 => x"4bc04a71",
   764 => x"c0029a72",
   765 => x"a2da87e0",
   766 => x"4b699f49",
   767 => x"bff0fec2",
   768 => x"d487cf02",
   769 => x"699f49a2",
   770 => x"ffc04c49",
   771 => x"34d09cff",
   772 => x"4cc087c2",
   773 => x"9b73b374",
   774 => x"4a87df02",
   775 => x"fec28ac2",
   776 => x"9249bfe8",
   777 => x"bfccc3c3",
   778 => x"c3807248",
   779 => x"7158ecc3",
   780 => x"c230c448",
   781 => x"c058f8fe",
   782 => x"c3c387e9",
   783 => x"c34bbfd0",
   784 => x"c348e8c3",
   785 => x"78bfd4c3",
   786 => x"bff0fec2",
   787 => x"c287c902",
   788 => x"49bfe8fe",
   789 => x"87c731c4",
   790 => x"bfd8c3c3",
   791 => x"c231c449",
   792 => x"c359f8fe",
   793 => x"265be8c3",
   794 => x"264b264c",
   795 => x"5b5e0e4f",
   796 => x"f00e5d5c",
   797 => x"59a6c886",
   798 => x"ffffffcf",
   799 => x"7ec04cf8",
   800 => x"d80266c4",
   801 => x"e4f6c287",
   802 => x"c278c048",
   803 => x"c348dcf6",
   804 => x"78bfe8c3",
   805 => x"48e0f6c2",
   806 => x"bfe4c3c3",
   807 => x"c5ffc278",
   808 => x"c250c048",
   809 => x"49bff4fe",
   810 => x"bfe4f6c2",
   811 => x"03aa714a",
   812 => x"7287ccc4",
   813 => x"0599cf49",
   814 => x"c087eac0",
   815 => x"c248e8f9",
   816 => x"78bfdcf6",
   817 => x"1ee8f6c2",
   818 => x"bfdcf6c2",
   819 => x"dcf6c249",
   820 => x"78a1c148",
   821 => x"fddfff71",
   822 => x"c086c487",
   823 => x"c248e4f9",
   824 => x"cc78e8f6",
   825 => x"e4f9c087",
   826 => x"e0c048bf",
   827 => x"e8f9c080",
   828 => x"e4f6c258",
   829 => x"80c148bf",
   830 => x"58e8f6c2",
   831 => x"000e6427",
   832 => x"bf97bf00",
   833 => x"c2029d4d",
   834 => x"e5c387e5",
   835 => x"dec202ad",
   836 => x"e4f9c087",
   837 => x"a3cb4bbf",
   838 => x"cf4c1149",
   839 => x"d2c105ac",
   840 => x"df497587",
   841 => x"cd89c199",
   842 => x"f8fec291",
   843 => x"4aa3c181",
   844 => x"a3c35112",
   845 => x"c551124a",
   846 => x"51124aa3",
   847 => x"124aa3c7",
   848 => x"4aa3c951",
   849 => x"a3ce5112",
   850 => x"d051124a",
   851 => x"51124aa3",
   852 => x"124aa3d2",
   853 => x"4aa3d451",
   854 => x"a3d65112",
   855 => x"d851124a",
   856 => x"51124aa3",
   857 => x"124aa3dc",
   858 => x"4aa3de51",
   859 => x"7ec15112",
   860 => x"7487fcc0",
   861 => x"0599c849",
   862 => x"7487edc0",
   863 => x"0599d049",
   864 => x"e0c087d3",
   865 => x"ccc00266",
   866 => x"c0497387",
   867 => x"700f66e0",
   868 => x"d3c00298",
   869 => x"c0056e87",
   870 => x"fec287c6",
   871 => x"50c048f8",
   872 => x"bfe4f9c0",
   873 => x"87ebc248",
   874 => x"48c5ffc2",
   875 => x"c27e50c0",
   876 => x"49bff4fe",
   877 => x"bfe4f6c2",
   878 => x"04aa714a",
   879 => x"cf87f4fb",
   880 => x"f8ffffff",
   881 => x"e8c3c34c",
   882 => x"c8c005bf",
   883 => x"f0fec287",
   884 => x"fcc102bf",
   885 => x"e0f6c287",
   886 => x"c4eb49bf",
   887 => x"e4f6c287",
   888 => x"48a6c458",
   889 => x"bfe0f6c2",
   890 => x"f0fec278",
   891 => x"dbc002bf",
   892 => x"4966c487",
   893 => x"a9749974",
   894 => x"87c8c002",
   895 => x"c048a6c8",
   896 => x"87e7c078",
   897 => x"c148a6c8",
   898 => x"87dfc078",
   899 => x"cf4966c4",
   900 => x"a999f8ff",
   901 => x"87c8c002",
   902 => x"c048a6cc",
   903 => x"87c5c078",
   904 => x"c148a6cc",
   905 => x"48a6c878",
   906 => x"c87866cc",
   907 => x"e0c00566",
   908 => x"4966c487",
   909 => x"fec289c2",
   910 => x"914abfe8",
   911 => x"bfccc3c3",
   912 => x"dcf6c24a",
   913 => x"78a17248",
   914 => x"48e4f6c2",
   915 => x"d2f978c0",
   916 => x"cf48c087",
   917 => x"f8ffffff",
   918 => x"268ef04c",
   919 => x"264c264d",
   920 => x"004f264b",
   921 => x"00000000",
   922 => x"ffffffff",
   923 => x"48d0ff1e",
   924 => x"2678e0c0",
   925 => x"e9c11e4f",
   926 => x"497087f7",
   927 => x"87c60299",
   928 => x"05a9fbc0",
   929 => x"487187f0",
   930 => x"5e0e4f26",
   931 => x"710e5c5b",
   932 => x"c14cc04b",
   933 => x"7087dae9",
   934 => x"c0029949",
   935 => x"ecc087fa",
   936 => x"f3c002a9",
   937 => x"a9fbc087",
   938 => x"87ecc002",
   939 => x"acb766cc",
   940 => x"d087c703",
   941 => x"87c20266",
   942 => x"99715371",
   943 => x"c187c202",
   944 => x"ece8c184",
   945 => x"99497087",
   946 => x"c087cd02",
   947 => x"c702a9ec",
   948 => x"a9fbc087",
   949 => x"87d4ff05",
   950 => x"c30266d0",
   951 => x"7b97c087",
   952 => x"05a9fbc0",
   953 => x"4a7487c7",
   954 => x"c28a0ac0",
   955 => x"724a7487",
   956 => x"264c2648",
   957 => x"1e4f264b",
   958 => x"87f5e7c1",
   959 => x"c04a4970",
   960 => x"c904aaf0",
   961 => x"aaf9c087",
   962 => x"c087c301",
   963 => x"c1c18af0",
   964 => x"87c904aa",
   965 => x"01aadac1",
   966 => x"f7c087c3",
   967 => x"2648728a",
   968 => x"5b5e0e4f",
   969 => x"f80e5d5c",
   970 => x"c04c7186",
   971 => x"e3e7c17e",
   972 => x"c04bc087",
   973 => x"bf97c4ff",
   974 => x"04a9c049",
   975 => x"f4fc87cf",
   976 => x"c083c187",
   977 => x"bf97c4ff",
   978 => x"f106ab49",
   979 => x"c4ffc087",
   980 => x"d002bf97",
   981 => x"d8e6c187",
   982 => x"99497087",
   983 => x"c087c602",
   984 => x"f005a9ec",
   985 => x"c14bc087",
   986 => x"7087c6e6",
   987 => x"c0e6c14d",
   988 => x"58a6c887",
   989 => x"87f9e5c1",
   990 => x"83c14a70",
   991 => x"9749a4c8",
   992 => x"05ad4969",
   993 => x"a4c987da",
   994 => x"49699749",
   995 => x"05a966c4",
   996 => x"a4ca87ce",
   997 => x"49699749",
   998 => x"87c405aa",
   999 => x"87d07ec1",
  1000 => x"02adecc0",
  1001 => x"fbc087c6",
  1002 => x"87c405ad",
  1003 => x"7ec14bc0",
  1004 => x"f2fe026e",
  1005 => x"87f4fa87",
  1006 => x"8ef84873",
  1007 => x"4c264d26",
  1008 => x"4f264b26",
  1009 => x"1e731e00",
  1010 => x"c84bd4ff",
  1011 => x"d0ff4a66",
  1012 => x"78c5c848",
  1013 => x"c148d4ff",
  1014 => x"7b1178d4",
  1015 => x"f9058ac1",
  1016 => x"48d0ff87",
  1017 => x"4b2678c4",
  1018 => x"5e0e4f26",
  1019 => x"0e5d5c5b",
  1020 => x"7e7186f8",
  1021 => x"c3c31e6e",
  1022 => x"dbe449fc",
  1023 => x"7086c487",
  1024 => x"e4c40298",
  1025 => x"e4e8c187",
  1026 => x"496e4cbf",
  1027 => x"c887d2fc",
  1028 => x"987058a6",
  1029 => x"c487c505",
  1030 => x"78c148a6",
  1031 => x"c548d0ff",
  1032 => x"48d4ff78",
  1033 => x"c478d5c1",
  1034 => x"89c14966",
  1035 => x"e8c131c6",
  1036 => x"4abf97dc",
  1037 => x"ffb07148",
  1038 => x"ff7808d4",
  1039 => x"78c448d0",
  1040 => x"97f8c3c3",
  1041 => x"99d049bf",
  1042 => x"c587dd02",
  1043 => x"48d4ff78",
  1044 => x"c078d6c1",
  1045 => x"48d4ff4a",
  1046 => x"c178ffc3",
  1047 => x"aae0c082",
  1048 => x"ff87f204",
  1049 => x"78c448d0",
  1050 => x"c348d4ff",
  1051 => x"d0ff78ff",
  1052 => x"ff78c548",
  1053 => x"d3c148d4",
  1054 => x"ff78c178",
  1055 => x"78c448d0",
  1056 => x"06acb7c0",
  1057 => x"c387cbc2",
  1058 => x"4bbfc4c4",
  1059 => x"737e748c",
  1060 => x"ddc1029b",
  1061 => x"4dc0c887",
  1062 => x"abb7c08b",
  1063 => x"c887c603",
  1064 => x"c04da3c0",
  1065 => x"f8c3c34b",
  1066 => x"d049bf97",
  1067 => x"87cf0299",
  1068 => x"c3c31ec0",
  1069 => x"d5e649fc",
  1070 => x"7086c487",
  1071 => x"c287d84c",
  1072 => x"c31ee8f6",
  1073 => x"e649fcc3",
  1074 => x"4c7087c4",
  1075 => x"f6c21e75",
  1076 => x"f0fb49e8",
  1077 => x"7486c887",
  1078 => x"87c5059c",
  1079 => x"cac148c0",
  1080 => x"c31ec187",
  1081 => x"e449fcc3",
  1082 => x"86c487d5",
  1083 => x"fe059b73",
  1084 => x"4c6e87e3",
  1085 => x"06acb7c0",
  1086 => x"c3c387d1",
  1087 => x"78c048fc",
  1088 => x"78c080d0",
  1089 => x"c4c380f4",
  1090 => x"c078bfc8",
  1091 => x"fd01acb7",
  1092 => x"d0ff87f5",
  1093 => x"ff78c548",
  1094 => x"d3c148d4",
  1095 => x"ff78c078",
  1096 => x"78c448d0",
  1097 => x"c2c048c1",
  1098 => x"f848c087",
  1099 => x"264d268e",
  1100 => x"264b264c",
  1101 => x"5b5e0e4f",
  1102 => x"fc0e5d5c",
  1103 => x"c04d7186",
  1104 => x"04ad4c4b",
  1105 => x"c087e8c0",
  1106 => x"741ee1fc",
  1107 => x"87c4029c",
  1108 => x"87c24ac0",
  1109 => x"49724ac1",
  1110 => x"c487d2ec",
  1111 => x"c17e7086",
  1112 => x"c2056e83",
  1113 => x"c14b7587",
  1114 => x"06ab7584",
  1115 => x"6e87d8ff",
  1116 => x"268efc48",
  1117 => x"264c264d",
  1118 => x"0e4f264b",
  1119 => x"5d5c5b5e",
  1120 => x"7186fc0e",
  1121 => x"91de494c",
  1122 => x"4ddcc5c3",
  1123 => x"6d978571",
  1124 => x"87ddc102",
  1125 => x"bfccc5c3",
  1126 => x"71817449",
  1127 => x"7087d6fe",
  1128 => x"0298487e",
  1129 => x"c387f3c0",
  1130 => x"704bd0c5",
  1131 => x"fe49cb4a",
  1132 => x"7487cdfd",
  1133 => x"c193cc4b",
  1134 => x"c483e8e8",
  1135 => x"fcc7c183",
  1136 => x"c149747b",
  1137 => x"7587d5c4",
  1138 => x"e0e8c17b",
  1139 => x"1e49bf97",
  1140 => x"49d0c5c3",
  1141 => x"87e9e5c1",
  1142 => x"497486c4",
  1143 => x"87fcc3c1",
  1144 => x"c5c149c0",
  1145 => x"c3c387d7",
  1146 => x"50c048f4",
  1147 => x"c7e0c049",
  1148 => x"268efc87",
  1149 => x"264c264d",
  1150 => x"004f264b",
  1151 => x"64616f4c",
  1152 => x"2e676e69",
  1153 => x"00002e2e",
  1154 => x"61422080",
  1155 => x"00006b63",
  1156 => x"64616f4c",
  1157 => x"202e2a20",
  1158 => x"00000000",
  1159 => x"0000203a",
  1160 => x"61422080",
  1161 => x"00006b63",
  1162 => x"78452080",
  1163 => x"00007469",
  1164 => x"49204453",
  1165 => x"2e74696e",
  1166 => x"0000002e",
  1167 => x"00004b4f",
  1168 => x"544f4f42",
  1169 => x"20202020",
  1170 => x"004d4f52",
  1171 => x"711e731e",
  1172 => x"c5c3494b",
  1173 => x"7181bfcc",
  1174 => x"7087dafb",
  1175 => x"c4029a4a",
  1176 => x"c2e64987",
  1177 => x"ccc5c387",
  1178 => x"7378c048",
  1179 => x"87fac149",
  1180 => x"4f264b26",
  1181 => x"711e731e",
  1182 => x"4aa3c44b",
  1183 => x"87d0c102",
  1184 => x"dc028ac1",
  1185 => x"c0028a87",
  1186 => x"058a87f2",
  1187 => x"c387d3c1",
  1188 => x"02bfccc5",
  1189 => x"4887cbc1",
  1190 => x"c5c388c1",
  1191 => x"c1c158d0",
  1192 => x"ccc5c387",
  1193 => x"89c649bf",
  1194 => x"59d0c5c3",
  1195 => x"03a9b7c0",
  1196 => x"c387efc0",
  1197 => x"c048ccc5",
  1198 => x"87e6c078",
  1199 => x"bfc8c5c3",
  1200 => x"c387df02",
  1201 => x"48bfccc5",
  1202 => x"c5c380c1",
  1203 => x"87d258d0",
  1204 => x"bfc8c5c3",
  1205 => x"c387cb02",
  1206 => x"48bfccc5",
  1207 => x"c5c380c6",
  1208 => x"497358d0",
  1209 => x"4b2687c4",
  1210 => x"5e0e4f26",
  1211 => x"0e5d5c5b",
  1212 => x"a6d086f0",
  1213 => x"e8f6c259",
  1214 => x"c34cc04d",
  1215 => x"c148c8c5",
  1216 => x"48a6c478",
  1217 => x"7e7578c0",
  1218 => x"bfccc5c3",
  1219 => x"06a8c048",
  1220 => x"7587fac0",
  1221 => x"e8f6c27e",
  1222 => x"c0029848",
  1223 => x"fcc087ef",
  1224 => x"66c81ee1",
  1225 => x"c087c402",
  1226 => x"c187c24d",
  1227 => x"e449754d",
  1228 => x"86c487fb",
  1229 => x"84c17e70",
  1230 => x"c14866c4",
  1231 => x"58a6c880",
  1232 => x"bfccc5c3",
  1233 => x"87c503ac",
  1234 => x"d1ff056e",
  1235 => x"c04d6e87",
  1236 => x"029d754c",
  1237 => x"c087e0c3",
  1238 => x"c81ee1fc",
  1239 => x"87c70266",
  1240 => x"c048a6cc",
  1241 => x"cc87c578",
  1242 => x"78c148a6",
  1243 => x"e34966cc",
  1244 => x"86c487fb",
  1245 => x"98487e70",
  1246 => x"87e8c202",
  1247 => x"9781cb49",
  1248 => x"99d04969",
  1249 => x"87d6c102",
  1250 => x"4accc9c1",
  1251 => x"91cc4974",
  1252 => x"81e8e8c1",
  1253 => x"81c87972",
  1254 => x"7451ffc3",
  1255 => x"c391de49",
  1256 => x"714ddcc5",
  1257 => x"97c1c285",
  1258 => x"49a5c17d",
  1259 => x"c251e0c0",
  1260 => x"bf97f8fe",
  1261 => x"c187d202",
  1262 => x"4ba5c284",
  1263 => x"4af8fec2",
  1264 => x"f4fe49db",
  1265 => x"dbc187fa",
  1266 => x"49a5cd87",
  1267 => x"84c151c0",
  1268 => x"6e4ba5c2",
  1269 => x"fe49cb4a",
  1270 => x"c187e5f4",
  1271 => x"c5c187c6",
  1272 => x"49744afb",
  1273 => x"e8c191cc",
  1274 => x"797281e8",
  1275 => x"97f8fec2",
  1276 => x"87d802bf",
  1277 => x"91de4974",
  1278 => x"c5c384c1",
  1279 => x"83714bdc",
  1280 => x"4af8fec2",
  1281 => x"f3fe49dd",
  1282 => x"87d887f6",
  1283 => x"93de4b74",
  1284 => x"83dcc5c3",
  1285 => x"c049a3cb",
  1286 => x"7384c151",
  1287 => x"49cb4a6e",
  1288 => x"87dcf3fe",
  1289 => x"c14866c4",
  1290 => x"58a6c880",
  1291 => x"c003acc7",
  1292 => x"056e87c5",
  1293 => x"c787e0fc",
  1294 => x"e6c003ac",
  1295 => x"c8c5c387",
  1296 => x"c178c048",
  1297 => x"744afbc5",
  1298 => x"c191cc49",
  1299 => x"7281e8e8",
  1300 => x"de497479",
  1301 => x"dcc5c391",
  1302 => x"c151c081",
  1303 => x"04acc784",
  1304 => x"c187daff",
  1305 => x"c048c4ea",
  1306 => x"c180f750",
  1307 => x"c140d1d3",
  1308 => x"c878c8c8",
  1309 => x"f4c9c180",
  1310 => x"4966cc78",
  1311 => x"87dcf9c0",
  1312 => x"4d268ef0",
  1313 => x"4b264c26",
  1314 => x"731e4f26",
  1315 => x"494b711e",
  1316 => x"e8c191cc",
  1317 => x"a1c881e8",
  1318 => x"dce8c14a",
  1319 => x"c9501248",
  1320 => x"ffc04aa1",
  1321 => x"501248c4",
  1322 => x"e8c181ca",
  1323 => x"501148e0",
  1324 => x"97e0e8c1",
  1325 => x"c01e49bf",
  1326 => x"c4dac149",
  1327 => x"f8497387",
  1328 => x"8efc87e8",
  1329 => x"4f264b26",
  1330 => x"c049c01e",
  1331 => x"2687eef9",
  1332 => x"4a711e4f",
  1333 => x"c191cc49",
  1334 => x"c881e8e8",
  1335 => x"f4c3c381",
  1336 => x"c0501148",
  1337 => x"fe49a2f0",
  1338 => x"c087e1ee",
  1339 => x"87c8d449",
  1340 => x"5e0e4f26",
  1341 => x"0e5d5c5b",
  1342 => x"4d7186f4",
  1343 => x"c191cc49",
  1344 => x"c881e8e8",
  1345 => x"a1ca4aa1",
  1346 => x"48a6c47e",
  1347 => x"bff0c3c3",
  1348 => x"bf976e78",
  1349 => x"4c66c44b",
  1350 => x"48122c73",
  1351 => x"7058a6cc",
  1352 => x"c984c19c",
  1353 => x"49699781",
  1354 => x"c204acb7",
  1355 => x"6e4cc087",
  1356 => x"c84abf97",
  1357 => x"31724966",
  1358 => x"66c4b9ff",
  1359 => x"72487499",
  1360 => x"b14a7030",
  1361 => x"59f4c3c3",
  1362 => x"f8cdc171",
  1363 => x"c31ec787",
  1364 => x"1ebfc4c5",
  1365 => x"1ee8e8c1",
  1366 => x"97f4c3c3",
  1367 => x"e2c149bf",
  1368 => x"c0497587",
  1369 => x"e887f5f5",
  1370 => x"264d268e",
  1371 => x"264b264c",
  1372 => x"1e731e4f",
  1373 => x"a3c24b71",
  1374 => x"87d6024a",
  1375 => x"c0058ac1",
  1376 => x"c5c387e2",
  1377 => x"db02bfc4",
  1378 => x"88c14887",
  1379 => x"58c8c5c3",
  1380 => x"c5c387d2",
  1381 => x"cb02bfc8",
  1382 => x"c4c5c387",
  1383 => x"80c148bf",
  1384 => x"58c8c5c3",
  1385 => x"c5c31ec7",
  1386 => x"c11ebfc4",
  1387 => x"c31ee8e8",
  1388 => x"bf97f4c3",
  1389 => x"7387cc49",
  1390 => x"dff4c049",
  1391 => x"268ef487",
  1392 => x"0e4f264b",
  1393 => x"5d5c5b5e",
  1394 => x"86ccff0e",
  1395 => x"59a6e8c0",
  1396 => x"c048a6cc",
  1397 => x"c080c478",
  1398 => x"c080c478",
  1399 => x"c180c478",
  1400 => x"c47866c8",
  1401 => x"c478c180",
  1402 => x"c378c180",
  1403 => x"c148c8c5",
  1404 => x"dfccc178",
  1405 => x"87fde187",
  1406 => x"87f5cbc1",
  1407 => x"fbc04d70",
  1408 => x"f2c102ad",
  1409 => x"66e4c087",
  1410 => x"87e7c105",
  1411 => x"4a66c4c1",
  1412 => x"7e6a82c4",
  1413 => x"48d0c8c1",
  1414 => x"4120496e",
  1415 => x"51104120",
  1416 => x"4866c4c1",
  1417 => x"78cad2c1",
  1418 => x"81c7496a",
  1419 => x"c4c15175",
  1420 => x"81c84966",
  1421 => x"a6dc51c1",
  1422 => x"c178c248",
  1423 => x"c94966c4",
  1424 => x"c151c081",
  1425 => x"ca4966c4",
  1426 => x"c151c081",
  1427 => x"6a1ed81e",
  1428 => x"e081c849",
  1429 => x"86c887f4",
  1430 => x"4866c8c1",
  1431 => x"c701a8c0",
  1432 => x"48a6d487",
  1433 => x"87cf78c1",
  1434 => x"4866c8c1",
  1435 => x"a6dc88c1",
  1436 => x"ff87c458",
  1437 => x"7587fedf",
  1438 => x"f3cb029d",
  1439 => x"4866d487",
  1440 => x"a866ccc1",
  1441 => x"87e8cb03",
  1442 => x"c9c17ec0",
  1443 => x"4d7087e3",
  1444 => x"88c6c148",
  1445 => x"7058a6c8",
  1446 => x"d6c10298",
  1447 => x"88c94887",
  1448 => x"7058a6c8",
  1449 => x"d9c50298",
  1450 => x"88c14887",
  1451 => x"7058a6c8",
  1452 => x"f8c20298",
  1453 => x"88c34887",
  1454 => x"7058a6c8",
  1455 => x"87cf0298",
  1456 => x"c888c148",
  1457 => x"987058a6",
  1458 => x"87f6c402",
  1459 => x"c087c0ca",
  1460 => x"c8c17ef0",
  1461 => x"4d7087db",
  1462 => x"02adecc0",
  1463 => x"7e7587c2",
  1464 => x"02adecc0",
  1465 => x"c8c187cd",
  1466 => x"4d7087c7",
  1467 => x"05adecc0",
  1468 => x"c087f3ff",
  1469 => x"c10566e4",
  1470 => x"ecc087ea",
  1471 => x"87c402ad",
  1472 => x"87edc7c1",
  1473 => x"1eca1ec0",
  1474 => x"cc4b66dc",
  1475 => x"66ccc193",
  1476 => x"4ca3c483",
  1477 => x"ddff496c",
  1478 => x"1ec187f0",
  1479 => x"496c1ede",
  1480 => x"87e6ddff",
  1481 => x"d2c186d0",
  1482 => x"a3c87bca",
  1483 => x"5166dc49",
  1484 => x"c049a3c9",
  1485 => x"ca5166e0",
  1486 => x"516e49a3",
  1487 => x"c14866dc",
  1488 => x"a6e0c080",
  1489 => x"4866d458",
  1490 => x"04a866d8",
  1491 => x"66d487cb",
  1492 => x"d880c148",
  1493 => x"fcc758a6",
  1494 => x"4866d887",
  1495 => x"a6dc88c1",
  1496 => x"87f1c758",
  1497 => x"87cddcff",
  1498 => x"e8c74d70",
  1499 => x"c6deff87",
  1500 => x"58a6d087",
  1501 => x"06a866d0",
  1502 => x"d087c6c0",
  1503 => x"66cc48a6",
  1504 => x"f2ddff78",
  1505 => x"a8ecc087",
  1506 => x"87f6c105",
  1507 => x"0566e4c0",
  1508 => x"d487e6c1",
  1509 => x"91cc4966",
  1510 => x"8166c4c1",
  1511 => x"6a4aa1c4",
  1512 => x"4aa1c84c",
  1513 => x"c15266cc",
  1514 => x"c179d1d3",
  1515 => x"7087c2c5",
  1516 => x"db029d4d",
  1517 => x"adfbc087",
  1518 => x"87d4c002",
  1519 => x"c4c15475",
  1520 => x"4d7087ef",
  1521 => x"c7c0029d",
  1522 => x"adfbc087",
  1523 => x"87ecff05",
  1524 => x"c254e0c0",
  1525 => x"97c054c1",
  1526 => x"4866d47c",
  1527 => x"04a866d8",
  1528 => x"d487cbc0",
  1529 => x"80c14866",
  1530 => x"c558a6d8",
  1531 => x"66d887e7",
  1532 => x"dc88c148",
  1533 => x"dcc558a6",
  1534 => x"f8d9ff87",
  1535 => x"c54d7087",
  1536 => x"66cc87d3",
  1537 => x"66e4c048",
  1538 => x"f4c405a8",
  1539 => x"a6e8c087",
  1540 => x"ff78c048",
  1541 => x"7087e0db",
  1542 => x"dadbff7e",
  1543 => x"a6f0c087",
  1544 => x"a8ecc058",
  1545 => x"87c7c005",
  1546 => x"786e48a6",
  1547 => x"c187c4c0",
  1548 => x"d487fec2",
  1549 => x"91cc4966",
  1550 => x"4866c4c1",
  1551 => x"a6c88071",
  1552 => x"4a66c458",
  1553 => x"66c482c8",
  1554 => x"6e81ca49",
  1555 => x"66ecc051",
  1556 => x"6e81c149",
  1557 => x"7148c189",
  1558 => x"c1497030",
  1559 => x"7a977189",
  1560 => x"bff0c3c3",
  1561 => x"97296e49",
  1562 => x"71484a6a",
  1563 => x"a6f4c098",
  1564 => x"4866c458",
  1565 => x"a6cc80c4",
  1566 => x"bf66c858",
  1567 => x"66e4c04c",
  1568 => x"a866cc48",
  1569 => x"87c5c002",
  1570 => x"c2c07ec0",
  1571 => x"6e7ec187",
  1572 => x"1ee0c01e",
  1573 => x"d7ff4974",
  1574 => x"86c887f0",
  1575 => x"b7c04d70",
  1576 => x"d4c106ad",
  1577 => x"c8847587",
  1578 => x"c049bf66",
  1579 => x"897481e0",
  1580 => x"dcc8c14b",
  1581 => x"e1fe714a",
  1582 => x"84c287c6",
  1583 => x"e8c07e74",
  1584 => x"80c14866",
  1585 => x"58a6ecc0",
  1586 => x"4966f0c0",
  1587 => x"a97081c1",
  1588 => x"87c5c002",
  1589 => x"c2c04cc0",
  1590 => x"744cc187",
  1591 => x"bf66cc1e",
  1592 => x"81e0c049",
  1593 => x"718966c4",
  1594 => x"4966c81e",
  1595 => x"87dad6ff",
  1596 => x"b7c086c8",
  1597 => x"c5ff01a8",
  1598 => x"66e8c087",
  1599 => x"87d3c002",
  1600 => x"c94966c4",
  1601 => x"66e8c081",
  1602 => x"4866c451",
  1603 => x"78f2d3c1",
  1604 => x"c487cec0",
  1605 => x"81c94966",
  1606 => x"66c451c2",
  1607 => x"e3ebc248",
  1608 => x"4866d478",
  1609 => x"04a866d8",
  1610 => x"d487cbc0",
  1611 => x"80c14866",
  1612 => x"c058a6d8",
  1613 => x"66d887d1",
  1614 => x"dc88c148",
  1615 => x"c6c058a6",
  1616 => x"f0d4ff87",
  1617 => x"cc4d7087",
  1618 => x"78c048a6",
  1619 => x"ff87c6c0",
  1620 => x"7087e2d4",
  1621 => x"66e0c04d",
  1622 => x"c080c148",
  1623 => x"7558a6e4",
  1624 => x"cbc0029d",
  1625 => x"4866d487",
  1626 => x"a866ccc1",
  1627 => x"87d8f404",
  1628 => x"c74866d4",
  1629 => x"e1c003a8",
  1630 => x"4c66d487",
  1631 => x"48c8c5c3",
  1632 => x"497478c0",
  1633 => x"c4c191cc",
  1634 => x"a1c48166",
  1635 => x"c04a6a4a",
  1636 => x"84c17952",
  1637 => x"ff04acc7",
  1638 => x"e4c087e2",
  1639 => x"e2c00266",
  1640 => x"66c4c187",
  1641 => x"81d4c149",
  1642 => x"4a66c4c1",
  1643 => x"c082dcc1",
  1644 => x"d1d3c152",
  1645 => x"66c4c179",
  1646 => x"81d8c149",
  1647 => x"79e0c8c1",
  1648 => x"c187d6c0",
  1649 => x"c14966c4",
  1650 => x"c4c181d4",
  1651 => x"d8c14a66",
  1652 => x"e8c8c182",
  1653 => x"c8d3c17a",
  1654 => x"f1d5c179",
  1655 => x"66c4c14a",
  1656 => x"81e0c149",
  1657 => x"d2ff7972",
  1658 => x"66d087c2",
  1659 => x"8eccff48",
  1660 => x"4c264d26",
  1661 => x"4f264b26",
  1662 => x"c31ec71e",
  1663 => x"1ebfc4c5",
  1664 => x"1ee8e8c1",
  1665 => x"97f4c3c3",
  1666 => x"f6ee49bf",
  1667 => x"e8e8c187",
  1668 => x"d5e4c049",
  1669 => x"268ef487",
  1670 => x"0000004f",
  1671 => x"00000000",
  1672 => x"00000000",
  1673 => x"00000001",
  1674 => x"0000117b",
  1675 => x"0000315c",
  1676 => x"00000000",
  1677 => x"0000117b",
  1678 => x"0000317a",
  1679 => x"00000000",
  1680 => x"0000117b",
  1681 => x"00003198",
  1682 => x"00000000",
  1683 => x"0000117b",
  1684 => x"000031b6",
  1685 => x"00000000",
  1686 => x"0000117b",
  1687 => x"000031d4",
  1688 => x"00000000",
  1689 => x"0000117b",
  1690 => x"000031f2",
  1691 => x"00000000",
  1692 => x"0000117b",
  1693 => x"00003210",
  1694 => x"00000000",
  1695 => x"000014d1",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00001274",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00001240",
  1702 => x"db86fc1e",
  1703 => x"fc7e7087",
  1704 => x"1e4f268e",
  1705 => x"c048f0fe",
  1706 => x"7909cd78",
  1707 => x"1e4f2609",
  1708 => x"49d8eac1",
  1709 => x"4f2687ed",
  1710 => x"bff0fe1e",
  1711 => x"1e4f2648",
  1712 => x"c148f0fe",
  1713 => x"1e4f2678",
  1714 => x"c048f0fe",
  1715 => x"1e4f2678",
  1716 => x"97c04a71",
  1717 => x"49a2c17a",
  1718 => x"a2ca51c0",
  1719 => x"cb51c049",
  1720 => x"51c049a2",
  1721 => x"5e0e4f26",
  1722 => x"f00e5c5b",
  1723 => x"ca4c7186",
  1724 => x"699749a4",
  1725 => x"4ba4cb7e",
  1726 => x"c8486b97",
  1727 => x"80c158a6",
  1728 => x"c758a6cc",
  1729 => x"58a6d098",
  1730 => x"66cc486e",
  1731 => x"87db05a8",
  1732 => x"977e6997",
  1733 => x"a6c8486b",
  1734 => x"cc80c158",
  1735 => x"98c758a6",
  1736 => x"6e58a6d0",
  1737 => x"a866cc48",
  1738 => x"fe87e502",
  1739 => x"a4cc87d9",
  1740 => x"496b974a",
  1741 => x"dc49a172",
  1742 => x"6b975166",
  1743 => x"c1486e7e",
  1744 => x"58a6c880",
  1745 => x"a6cc98c7",
  1746 => x"7b977058",
  1747 => x"fd87dec1",
  1748 => x"8ef087ed",
  1749 => x"4b264c26",
  1750 => x"5e0e4f26",
  1751 => x"0e5d5c5b",
  1752 => x"4d7186f4",
  1753 => x"c17e6d97",
  1754 => x"6c974ca5",
  1755 => x"58a6c848",
  1756 => x"66c4486e",
  1757 => x"87c505a8",
  1758 => x"e6c048ff",
  1759 => x"87c7fd87",
  1760 => x"9749a5c2",
  1761 => x"a3714b6c",
  1762 => x"4b6b974b",
  1763 => x"6e7e6c97",
  1764 => x"c880c148",
  1765 => x"98c758a6",
  1766 => x"7058a6cc",
  1767 => x"defc7c97",
  1768 => x"f4487387",
  1769 => x"264d268e",
  1770 => x"264b264c",
  1771 => x"5b5e0e4f",
  1772 => x"86f40e5c",
  1773 => x"e087d0fc",
  1774 => x"c0494cbf",
  1775 => x"0299c0e0",
  1776 => x"7487eac0",
  1777 => x"9affc34a",
  1778 => x"97c4c9c3",
  1779 => x"c9c349bf",
  1780 => x"517281c6",
  1781 => x"97c4c9c3",
  1782 => x"486e7ebf",
  1783 => x"a6c880c1",
  1784 => x"cc98c758",
  1785 => x"c9c358a6",
  1786 => x"66c848c4",
  1787 => x"d0497450",
  1788 => x"c10299c0",
  1789 => x"c9c387c0",
  1790 => x"7ebf97ce",
  1791 => x"97cfc9c3",
  1792 => x"a6c848bf",
  1793 => x"c4486e58",
  1794 => x"c002a866",
  1795 => x"c9c387e8",
  1796 => x"49bf97ce",
  1797 => x"81d0c9c3",
  1798 => x"08e04811",
  1799 => x"cec9c378",
  1800 => x"6e7ebf97",
  1801 => x"c880c148",
  1802 => x"98c758a6",
  1803 => x"c358a6cc",
  1804 => x"c848cec9",
  1805 => x"bfe45066",
  1806 => x"e0c0494b",
  1807 => x"c00299c0",
  1808 => x"4a7387ea",
  1809 => x"c39affc3",
  1810 => x"bf97d8c9",
  1811 => x"dac9c349",
  1812 => x"c3517281",
  1813 => x"bf97d8c9",
  1814 => x"c1486e7e",
  1815 => x"58a6c880",
  1816 => x"a6cc98c7",
  1817 => x"d8c9c358",
  1818 => x"5066c848",
  1819 => x"c0d04973",
  1820 => x"c0c10299",
  1821 => x"e2c9c387",
  1822 => x"c37ebf97",
  1823 => x"bf97e3c9",
  1824 => x"58a6c848",
  1825 => x"66c4486e",
  1826 => x"e8c002a8",
  1827 => x"e2c9c387",
  1828 => x"c349bf97",
  1829 => x"1181e4c9",
  1830 => x"7808e448",
  1831 => x"97e2c9c3",
  1832 => x"486e7ebf",
  1833 => x"a6c880c1",
  1834 => x"cc98c758",
  1835 => x"c9c358a6",
  1836 => x"66c848e2",
  1837 => x"87c0f850",
  1838 => x"c2f87e70",
  1839 => x"268ef487",
  1840 => x"264b264c",
  1841 => x"c9c31e4f",
  1842 => x"c2f849c4",
  1843 => x"d8c9c387",
  1844 => x"87fbf749",
  1845 => x"49edeec1",
  1846 => x"c387c8f7",
  1847 => x"4f2687f2",
  1848 => x"c31e731e",
  1849 => x"f949c4c9",
  1850 => x"4a7087f0",
  1851 => x"04aab7c0",
  1852 => x"c387ccc2",
  1853 => x"c905aaf0",
  1854 => x"c8f6c187",
  1855 => x"c178c148",
  1856 => x"e0c387ed",
  1857 => x"87c905aa",
  1858 => x"48ccf6c1",
  1859 => x"dec178c1",
  1860 => x"ccf6c187",
  1861 => x"87c602bf",
  1862 => x"4ba2c0c2",
  1863 => x"4b7287c2",
  1864 => x"bfc8f6c1",
  1865 => x"87e0c002",
  1866 => x"b7c44973",
  1867 => x"f6c19129",
  1868 => x"4a7381d0",
  1869 => x"92c29acf",
  1870 => x"307248c1",
  1871 => x"baff4a70",
  1872 => x"98694872",
  1873 => x"87db7970",
  1874 => x"b7c44973",
  1875 => x"f6c19129",
  1876 => x"4a7381d0",
  1877 => x"92c29acf",
  1878 => x"307248c3",
  1879 => x"69484a70",
  1880 => x"c17970b0",
  1881 => x"c048ccf6",
  1882 => x"c8f6c178",
  1883 => x"c378c048",
  1884 => x"f749c4c9",
  1885 => x"4a7087e4",
  1886 => x"03aab7c0",
  1887 => x"c087f4fd",
  1888 => x"264b2648",
  1889 => x"0000004f",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"00000000",
  1894 => x"00000000",
  1895 => x"00000000",
  1896 => x"00000000",
  1897 => x"00000000",
  1898 => x"00000000",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"724ac01e",
  1909 => x"c191c449",
  1910 => x"c081d0f6",
  1911 => x"d082c179",
  1912 => x"ee04aab7",
  1913 => x"0e4f2687",
  1914 => x"5d5c5b5e",
  1915 => x"f34d710e",
  1916 => x"4a7587d5",
  1917 => x"922ab7c4",
  1918 => x"82d0f6c1",
  1919 => x"9ccf4c75",
  1920 => x"496a94c2",
  1921 => x"c32b744b",
  1922 => x"7448c29b",
  1923 => x"ff4c7030",
  1924 => x"714874bc",
  1925 => x"f27a7098",
  1926 => x"487387e5",
  1927 => x"4c264d26",
  1928 => x"4f264b26",
  1929 => x"48d0ff1e",
  1930 => x"7178e1c8",
  1931 => x"08d4ff48",
  1932 => x"1e4f2678",
  1933 => x"c848d0ff",
  1934 => x"487178e1",
  1935 => x"7808d4ff",
  1936 => x"ff4866c4",
  1937 => x"267808d4",
  1938 => x"4a711e4f",
  1939 => x"1e4966c4",
  1940 => x"deff4972",
  1941 => x"48d0ff87",
  1942 => x"fc78e0c0",
  1943 => x"1e4f268e",
  1944 => x"4a711e73",
  1945 => x"abb7c24b",
  1946 => x"a387c803",
  1947 => x"ffc34a49",
  1948 => x"ce87c79a",
  1949 => x"c34a49a3",
  1950 => x"66c89aff",
  1951 => x"49721e49",
  1952 => x"fc87c6ff",
  1953 => x"264b268e",
  1954 => x"d0ff1e4f",
  1955 => x"78c9c848",
  1956 => x"d4ff4871",
  1957 => x"4f267808",
  1958 => x"494a711e",
  1959 => x"d0ff87eb",
  1960 => x"2678c848",
  1961 => x"1e731e4f",
  1962 => x"c9c34b71",
  1963 => x"c302bff8",
  1964 => x"87ebc287",
  1965 => x"c848d0ff",
  1966 => x"487378c9",
  1967 => x"ffb0e0c0",
  1968 => x"c37808d4",
  1969 => x"c048ecc9",
  1970 => x"0266c878",
  1971 => x"ffc387c5",
  1972 => x"c087c249",
  1973 => x"f4c9c349",
  1974 => x"0266cc59",
  1975 => x"d5c587c6",
  1976 => x"87c44ad5",
  1977 => x"4affffcf",
  1978 => x"5af8c9c3",
  1979 => x"48f8c9c3",
  1980 => x"4b2678c1",
  1981 => x"5e0e4f26",
  1982 => x"0e5d5c5b",
  1983 => x"c9c34d71",
  1984 => x"754bbff4",
  1985 => x"87cb029d",
  1986 => x"c191c849",
  1987 => x"714adcfa",
  1988 => x"c187c482",
  1989 => x"c04adcfe",
  1990 => x"7349124c",
  1991 => x"f0c9c399",
  1992 => x"b87148bf",
  1993 => x"7808d4ff",
  1994 => x"842bb7c1",
  1995 => x"04acb7c8",
  1996 => x"c9c387e7",
  1997 => x"c848bfec",
  1998 => x"f0c9c380",
  1999 => x"264d2658",
  2000 => x"264b264c",
  2001 => x"1e731e4f",
  2002 => x"4a134b71",
  2003 => x"87cb029a",
  2004 => x"e1fe4972",
  2005 => x"9a4a1387",
  2006 => x"2687f505",
  2007 => x"1e4f264b",
  2008 => x"bfecc9c3",
  2009 => x"ecc9c349",
  2010 => x"78a1c148",
  2011 => x"a9b7c0c4",
  2012 => x"ff87db03",
  2013 => x"c9c348d4",
  2014 => x"c378bff0",
  2015 => x"49bfecc9",
  2016 => x"48ecc9c3",
  2017 => x"c478a1c1",
  2018 => x"04a9b7c0",
  2019 => x"d0ff87e5",
  2020 => x"c378c848",
  2021 => x"c048f8c9",
  2022 => x"004f2678",
  2023 => x"00000000",
  2024 => x"00000000",
  2025 => x"5f000000",
  2026 => x"0000005f",
  2027 => x"00030300",
  2028 => x"00000303",
  2029 => x"147f7f14",
  2030 => x"00147f7f",
  2031 => x"6b2e2400",
  2032 => x"00123a6b",
  2033 => x"18366a4c",
  2034 => x"0032566c",
  2035 => x"594f7e30",
  2036 => x"40683a77",
  2037 => x"07040000",
  2038 => x"00000003",
  2039 => x"3e1c0000",
  2040 => x"00004163",
  2041 => x"63410000",
  2042 => x"00001c3e",
  2043 => x"1c3e2a08",
  2044 => x"082a3e1c",
  2045 => x"3e080800",
  2046 => x"0008083e",
  2047 => x"e0800000",
  2048 => x"00000060",
  2049 => x"08080800",
  2050 => x"00080808",
  2051 => x"60000000",
  2052 => x"00000060",
  2053 => x"18306040",
  2054 => x"0103060c",
  2055 => x"597f3e00",
  2056 => x"003e7f4d",
  2057 => x"7f060400",
  2058 => x"0000007f",
  2059 => x"71634200",
  2060 => x"00464f59",
  2061 => x"49632200",
  2062 => x"00367f49",
  2063 => x"13161c18",
  2064 => x"00107f7f",
  2065 => x"45672700",
  2066 => x"00397d45",
  2067 => x"4b7e3c00",
  2068 => x"00307949",
  2069 => x"71010100",
  2070 => x"00070f79",
  2071 => x"497f3600",
  2072 => x"00367f49",
  2073 => x"494f0600",
  2074 => x"001e3f69",
  2075 => x"66000000",
  2076 => x"00000066",
  2077 => x"e6800000",
  2078 => x"00000066",
  2079 => x"14080800",
  2080 => x"00222214",
  2081 => x"14141400",
  2082 => x"00141414",
  2083 => x"14222200",
  2084 => x"00080814",
  2085 => x"51030200",
  2086 => x"00060f59",
  2087 => x"5d417f3e",
  2088 => x"001e1f55",
  2089 => x"097f7e00",
  2090 => x"007e7f09",
  2091 => x"497f7f00",
  2092 => x"00367f49",
  2093 => x"633e1c00",
  2094 => x"00414141",
  2095 => x"417f7f00",
  2096 => x"001c3e63",
  2097 => x"497f7f00",
  2098 => x"00414149",
  2099 => x"097f7f00",
  2100 => x"00010109",
  2101 => x"417f3e00",
  2102 => x"007a7b49",
  2103 => x"087f7f00",
  2104 => x"007f7f08",
  2105 => x"7f410000",
  2106 => x"0000417f",
  2107 => x"40602000",
  2108 => x"003f7f40",
  2109 => x"1c087f7f",
  2110 => x"00416336",
  2111 => x"407f7f00",
  2112 => x"00404040",
  2113 => x"0c067f7f",
  2114 => x"007f7f06",
  2115 => x"0c067f7f",
  2116 => x"007f7f18",
  2117 => x"417f3e00",
  2118 => x"003e7f41",
  2119 => x"097f7f00",
  2120 => x"00060f09",
  2121 => x"61417f3e",
  2122 => x"00407e7f",
  2123 => x"097f7f00",
  2124 => x"00667f19",
  2125 => x"4d6f2600",
  2126 => x"00327b59",
  2127 => x"7f010100",
  2128 => x"0001017f",
  2129 => x"407f3f00",
  2130 => x"003f7f40",
  2131 => x"703f0f00",
  2132 => x"000f3f70",
  2133 => x"18307f7f",
  2134 => x"007f7f30",
  2135 => x"1c366341",
  2136 => x"4163361c",
  2137 => x"7c060301",
  2138 => x"0103067c",
  2139 => x"4d597161",
  2140 => x"00414347",
  2141 => x"7f7f0000",
  2142 => x"00004141",
  2143 => x"0c060301",
  2144 => x"40603018",
  2145 => x"41410000",
  2146 => x"00007f7f",
  2147 => x"03060c08",
  2148 => x"00080c06",
  2149 => x"80808080",
  2150 => x"00808080",
  2151 => x"03000000",
  2152 => x"00000407",
  2153 => x"54742000",
  2154 => x"00787c54",
  2155 => x"447f7f00",
  2156 => x"00387c44",
  2157 => x"447c3800",
  2158 => x"00004444",
  2159 => x"447c3800",
  2160 => x"007f7f44",
  2161 => x"547c3800",
  2162 => x"00185c54",
  2163 => x"7f7e0400",
  2164 => x"00000505",
  2165 => x"a4bc1800",
  2166 => x"007cfca4",
  2167 => x"047f7f00",
  2168 => x"00787c04",
  2169 => x"3d000000",
  2170 => x"0000407d",
  2171 => x"80808000",
  2172 => x"00007dfd",
  2173 => x"107f7f00",
  2174 => x"00446c38",
  2175 => x"3f000000",
  2176 => x"0000407f",
  2177 => x"180c7c7c",
  2178 => x"00787c0c",
  2179 => x"047c7c00",
  2180 => x"00787c04",
  2181 => x"447c3800",
  2182 => x"00387c44",
  2183 => x"24fcfc00",
  2184 => x"00183c24",
  2185 => x"243c1800",
  2186 => x"00fcfc24",
  2187 => x"047c7c00",
  2188 => x"00080c04",
  2189 => x"545c4800",
  2190 => x"00207454",
  2191 => x"7f3f0400",
  2192 => x"00004444",
  2193 => x"407c3c00",
  2194 => x"007c7c40",
  2195 => x"603c1c00",
  2196 => x"001c3c60",
  2197 => x"30607c3c",
  2198 => x"003c7c60",
  2199 => x"10386c44",
  2200 => x"00446c38",
  2201 => x"e0bc1c00",
  2202 => x"001c3c60",
  2203 => x"74644400",
  2204 => x"00444c5c",
  2205 => x"3e080800",
  2206 => x"00414177",
  2207 => x"7f000000",
  2208 => x"0000007f",
  2209 => x"77414100",
  2210 => x"0008083e",
  2211 => x"03010102",
  2212 => x"00010202",
  2213 => x"7f7f7f7f",
  2214 => x"007f7f7f",
  2215 => x"1c1c0808",
  2216 => x"7f7f3e3e",
  2217 => x"3e3e7f7f",
  2218 => x"08081c1c",
  2219 => x"7c181000",
  2220 => x"0010187c",
  2221 => x"7c301000",
  2222 => x"0010307c",
  2223 => x"60603010",
  2224 => x"00061e78",
  2225 => x"183c6642",
  2226 => x"0042663c",
  2227 => x"c26a3878",
  2228 => x"00386cc6",
  2229 => x"60000060",
  2230 => x"00600000",
  2231 => x"5c5b5e0e",
  2232 => x"86fc0e5d",
  2233 => x"cac37e71",
  2234 => x"c04cbfc0",
  2235 => x"c41ec04b",
  2236 => x"c402ab66",
  2237 => x"c24dc087",
  2238 => x"754dc187",
  2239 => x"ee49731e",
  2240 => x"86c887e3",
  2241 => x"ef49e0c0",
  2242 => x"a4c487ec",
  2243 => x"f0496a4a",
  2244 => x"caf187f3",
  2245 => x"c184cc87",
  2246 => x"abb7c883",
  2247 => x"87cdff04",
  2248 => x"4d268efc",
  2249 => x"4b264c26",
  2250 => x"711e4f26",
  2251 => x"c4cac34a",
  2252 => x"c4cac35a",
  2253 => x"4978c748",
  2254 => x"2687e1fe",
  2255 => x"1e731e4f",
  2256 => x"0bfc4b71",
  2257 => x"4a730b7b",
  2258 => x"c0c19ac1",
  2259 => x"c7ed49a2",
  2260 => x"d0dac287",
  2261 => x"264b265b",
  2262 => x"4a711e4f",
  2263 => x"721e66c4",
  2264 => x"87fbeb49",
  2265 => x"4f268efc",
  2266 => x"48d4ff1e",
  2267 => x"ff78ffc3",
  2268 => x"e1c048d0",
  2269 => x"48d4ff78",
  2270 => x"487178c1",
  2271 => x"d4ff30c4",
  2272 => x"d0ff7808",
  2273 => x"78e0c048",
  2274 => x"5e0e4f26",
  2275 => x"0e5d5c5b",
  2276 => x"7ec086f4",
  2277 => x"ec48a6c8",
  2278 => x"80fc78bf",
  2279 => x"bfc0cac3",
  2280 => x"c8cac378",
  2281 => x"bfe84cbf",
  2282 => x"ccdac24d",
  2283 => x"efe449bf",
  2284 => x"e849c787",
  2285 => x"497087f1",
  2286 => x"d00599c2",
  2287 => x"c4dac287",
  2288 => x"b9ff49bf",
  2289 => x"c19966c8",
  2290 => x"f9c10299",
  2291 => x"49e8cf87",
  2292 => x"7087fdca",
  2293 => x"e849c74b",
  2294 => x"987087cd",
  2295 => x"c887c905",
  2296 => x"99c14966",
  2297 => x"87fec002",
  2298 => x"ec48a6c8",
  2299 => x"efe378bf",
  2300 => x"ca497387",
  2301 => x"987087e6",
  2302 => x"c287d702",
  2303 => x"49bfc0da",
  2304 => x"dac2b9c1",
  2305 => x"fd7159c4",
  2306 => x"e8cf87de",
  2307 => x"87c0ca49",
  2308 => x"49c74b70",
  2309 => x"7087d0e7",
  2310 => x"cbff0598",
  2311 => x"4966c887",
  2312 => x"ff0599c1",
  2313 => x"dac287c2",
  2314 => x"c14abfcc",
  2315 => x"d0dac2ba",
  2316 => x"7a0afc5a",
  2317 => x"c19ac10a",
  2318 => x"e949a2c0",
  2319 => x"dac187da",
  2320 => x"87e3e649",
  2321 => x"dac27ec1",
  2322 => x"66c848c4",
  2323 => x"ccdac278",
  2324 => x"e9c005bf",
  2325 => x"c3497587",
  2326 => x"1e7199ff",
  2327 => x"f8fb49c0",
  2328 => x"c8497587",
  2329 => x"1e7129b7",
  2330 => x"ecfb49c1",
  2331 => x"c386c887",
  2332 => x"f2e549fd",
  2333 => x"49fac387",
  2334 => x"c787ece5",
  2335 => x"497587f4",
  2336 => x"c899ffc3",
  2337 => x"b5712db7",
  2338 => x"c0029d75",
  2339 => x"a6c887e4",
  2340 => x"bfc8ff48",
  2341 => x"4966c878",
  2342 => x"bfc8dac2",
  2343 => x"a9e0c289",
  2344 => x"87c4c003",
  2345 => x"87d04dc0",
  2346 => x"48c8dac2",
  2347 => x"c07866c8",
  2348 => x"dac287c6",
  2349 => x"78c048c8",
  2350 => x"99c84975",
  2351 => x"87cec005",
  2352 => x"e449f5c3",
  2353 => x"497087e1",
  2354 => x"c00299c2",
  2355 => x"cac387e7",
  2356 => x"c002bfc4",
  2357 => x"c14887ca",
  2358 => x"c8cac388",
  2359 => x"87d3c058",
  2360 => x"c14866c4",
  2361 => x"7e7080e0",
  2362 => x"c002bf6e",
  2363 => x"ff4b87c5",
  2364 => x"c10f7349",
  2365 => x"c449757e",
  2366 => x"cec00599",
  2367 => x"49f2c387",
  2368 => x"7087e4e3",
  2369 => x"0299c249",
  2370 => x"c387eac0",
  2371 => x"7ebfc4ca",
  2372 => x"a8b7c748",
  2373 => x"87cbc003",
  2374 => x"80c1486e",
  2375 => x"58c8cac3",
  2376 => x"c487d0c0",
  2377 => x"e0c14a66",
  2378 => x"c0026a82",
  2379 => x"fe4b87c5",
  2380 => x"c10f7349",
  2381 => x"49fdc37e",
  2382 => x"7087ece2",
  2383 => x"0299c249",
  2384 => x"c387e6c0",
  2385 => x"02bfc4ca",
  2386 => x"c387c9c0",
  2387 => x"c048c4ca",
  2388 => x"87d3c078",
  2389 => x"c14866c4",
  2390 => x"7e7080e0",
  2391 => x"c002bf6e",
  2392 => x"fd4b87c5",
  2393 => x"c10f7349",
  2394 => x"49fac37e",
  2395 => x"7087f8e1",
  2396 => x"0299c249",
  2397 => x"c387eac0",
  2398 => x"48bfc4ca",
  2399 => x"03a8b7c7",
  2400 => x"c387c9c0",
  2401 => x"c748c4ca",
  2402 => x"87d3c078",
  2403 => x"c14866c4",
  2404 => x"7e7080e0",
  2405 => x"c002bf6e",
  2406 => x"fc4b87c5",
  2407 => x"c10f7349",
  2408 => x"c348757e",
  2409 => x"a6cc98f0",
  2410 => x"05987058",
  2411 => x"c187cec0",
  2412 => x"f2e049da",
  2413 => x"c2497087",
  2414 => x"f9c10299",
  2415 => x"49e8cf87",
  2416 => x"7087cdc3",
  2417 => x"fcc9c34b",
  2418 => x"c350c048",
  2419 => x"bf97fcc9",
  2420 => x"87d2c105",
  2421 => x"c00566c8",
  2422 => x"dac187cc",
  2423 => x"87c7e049",
  2424 => x"c1029870",
  2425 => x"bfe887c0",
  2426 => x"ffc3494d",
  2427 => x"2db7c899",
  2428 => x"dbffb571",
  2429 => x"497387ea",
  2430 => x"7087e1c2",
  2431 => x"c6c00298",
  2432 => x"fcc9c387",
  2433 => x"c350c148",
  2434 => x"bf97fcc9",
  2435 => x"87d6c005",
  2436 => x"f0c34975",
  2437 => x"cdff0599",
  2438 => x"49dac187",
  2439 => x"87c7dfff",
  2440 => x"ff059870",
  2441 => x"cac387c0",
  2442 => x"4b49bfc4",
  2443 => x"66c493cc",
  2444 => x"714b6b83",
  2445 => x"9c740f73",
  2446 => x"87e9c002",
  2447 => x"e4c0026c",
  2448 => x"ff496c87",
  2449 => x"7087e0de",
  2450 => x"0299c149",
  2451 => x"c487cbc0",
  2452 => x"cac34ba4",
  2453 => x"6b49bfc4",
  2454 => x"84c80f4b",
  2455 => x"87c5c002",
  2456 => x"dcff056c",
  2457 => x"c0026e87",
  2458 => x"cac387c8",
  2459 => x"f149bfc4",
  2460 => x"8ef487ea",
  2461 => x"4c264d26",
  2462 => x"4f264b26",
  2463 => x"00000010",
  2464 => x"00000000",
  2465 => x"00000000",
  2466 => x"00000000",
  2467 => x"00000000",
  2468 => x"ff4a711e",
  2469 => x"7249bfc8",
  2470 => x"4f2648a1",
  2471 => x"bfc8ff1e",
  2472 => x"c0c0fe89",
  2473 => x"a9c0c0c0",
  2474 => x"c087c401",
  2475 => x"c187c24a",
  2476 => x"2648724a",
  2477 => x"5b5e0e4f",
  2478 => x"710e5d5c",
  2479 => x"4cd4ff4b",
  2480 => x"c04866d0",
  2481 => x"ff49d678",
  2482 => x"c387d9dd",
  2483 => x"496c7cff",
  2484 => x"7199ffc3",
  2485 => x"f0c3494d",
  2486 => x"a9e0c199",
  2487 => x"c387cb05",
  2488 => x"486c7cff",
  2489 => x"66d098c3",
  2490 => x"ffc37808",
  2491 => x"494a6c7c",
  2492 => x"ffc331c8",
  2493 => x"714a6c7c",
  2494 => x"c84972b2",
  2495 => x"7cffc331",
  2496 => x"b2714a6c",
  2497 => x"31c84972",
  2498 => x"6c7cffc3",
  2499 => x"ffb2714a",
  2500 => x"e0c048d0",
  2501 => x"029b7378",
  2502 => x"7b7287c2",
  2503 => x"4d264875",
  2504 => x"4b264c26",
  2505 => x"261e4f26",
  2506 => x"5b5e0e4f",
  2507 => x"86f80e5c",
  2508 => x"a6c81e76",
  2509 => x"87fdfd49",
  2510 => x"4b7086c4",
  2511 => x"a8c2486e",
  2512 => x"87fbc203",
  2513 => x"f0c34a73",
  2514 => x"aad0c19a",
  2515 => x"c187c702",
  2516 => x"c205aae0",
  2517 => x"497387e9",
  2518 => x"c30299c8",
  2519 => x"87c6ff87",
  2520 => x"9cc34c73",
  2521 => x"c105acc2",
  2522 => x"66c487c4",
  2523 => x"7131c949",
  2524 => x"4a66c41e",
  2525 => x"c392ccc1",
  2526 => x"7249ccca",
  2527 => x"cbcdfe81",
  2528 => x"ff49d887",
  2529 => x"c887ddda",
  2530 => x"f6c21ec0",
  2531 => x"e6fd49e8",
  2532 => x"d0ff87e1",
  2533 => x"78e0c048",
  2534 => x"1ee8f6c2",
  2535 => x"c14a66cc",
  2536 => x"cac392cc",
  2537 => x"817249cc",
  2538 => x"87e1cbfe",
  2539 => x"acc186cc",
  2540 => x"87cbc105",
  2541 => x"fd49eec0",
  2542 => x"c487d1e3",
  2543 => x"31c94966",
  2544 => x"66c41e71",
  2545 => x"92ccc14a",
  2546 => x"49cccac3",
  2547 => x"cbfe8172",
  2548 => x"f6c287fa",
  2549 => x"66c81ee8",
  2550 => x"92ccc14a",
  2551 => x"49cccac3",
  2552 => x"c9fe8172",
  2553 => x"49d787e8",
  2554 => x"87f8d8ff",
  2555 => x"c21ec0c8",
  2556 => x"fd49e8f6",
  2557 => x"cc87d9e4",
  2558 => x"48d0ff86",
  2559 => x"f878e0c0",
  2560 => x"264c268e",
  2561 => x"1e4f264b",
  2562 => x"b7c24a71",
  2563 => x"87ce03aa",
  2564 => x"ccc14972",
  2565 => x"cccac391",
  2566 => x"81c8c181",
  2567 => x"4f2679c0",
  2568 => x"5c5b5e0e",
  2569 => x"86fc0e5d",
  2570 => x"d4ff4a71",
  2571 => x"d44cc04b",
  2572 => x"b7c34d66",
  2573 => x"c2c201ad",
  2574 => x"029a7287",
  2575 => x"1e87ecc0",
  2576 => x"ccc14975",
  2577 => x"cccac391",
  2578 => x"c8807148",
  2579 => x"66c458a6",
  2580 => x"c3c3fe49",
  2581 => x"7086c487",
  2582 => x"87d40298",
  2583 => x"c8c1496e",
  2584 => x"6e79c181",
  2585 => x"6981c849",
  2586 => x"7587c54c",
  2587 => x"87d7fe49",
  2588 => x"c848d0ff",
  2589 => x"7bdd78e1",
  2590 => x"ffc34874",
  2591 => x"747b7098",
  2592 => x"29b7c849",
  2593 => x"ffc34871",
  2594 => x"747b7098",
  2595 => x"29b7d049",
  2596 => x"ffc34871",
  2597 => x"747b7098",
  2598 => x"28b7d848",
  2599 => x"7bc07b70",
  2600 => x"7b7b7b7b",
  2601 => x"7b7b7b7b",
  2602 => x"ff7b7b7b",
  2603 => x"e0c048d0",
  2604 => x"dc1e7578",
  2605 => x"d0d6ff49",
  2606 => x"fc86c487",
  2607 => x"264d268e",
  2608 => x"264b264c",
  2609 => x"d4ff1e4f",
  2610 => x"7affc34a",
  2611 => x"c548d0ff",
  2612 => x"717ac478",
  2613 => x"28b7d848",
  2614 => x"48717a70",
  2615 => x"7028b7d0",
  2616 => x"c848717a",
  2617 => x"7a7028b7",
  2618 => x"d0ff7a71",
  2619 => x"2678c448",
  2620 => x"4ac01e4f",
  2621 => x"bfe4ccc3",
  2622 => x"4987ca02",
  2623 => x"48e4ccc3",
  2624 => x"1178a1c1",
  2625 => x"059a724a",
  2626 => x"ccc387c6",
  2627 => x"78c048e4",
  2628 => x"4f264872",
  2629 => x"e4ccc31e",
  2630 => x"c0ebc248",
  2631 => x"4f2678bf",
  2632 => x"5c5b5e0e",
  2633 => x"ff4a710e",
  2634 => x"d4ff4cd0",
  2635 => x"c17cc54b",
  2636 => x"7bc37bd5",
  2637 => x"7cc57cc4",
  2638 => x"c17bd3c1",
  2639 => x"c87cc47b",
  2640 => x"d4c17cc5",
  2641 => x"b749c07b",
  2642 => x"87ca06aa",
  2643 => x"81c17bc0",
  2644 => x"04a9b772",
  2645 => x"7cc487f6",
  2646 => x"d3c17cc5",
  2647 => x"c47bc07b",
  2648 => x"264c267c",
  2649 => x"1e4f264b",
  2650 => x"4b711e73",
  2651 => x"fcc3c31e",
  2652 => x"e3fefd49",
  2653 => x"7086c487",
  2654 => x"e1c00298",
  2655 => x"c4c4c387",
  2656 => x"2aca4abf",
  2657 => x"028ac0c3",
  2658 => x"c0c187ce",
  2659 => x"87ce058a",
  2660 => x"48dce8c1",
  2661 => x"87c650c0",
  2662 => x"48dce8c1",
  2663 => x"4b2650c1",
  2664 => x"731e4f26",
  2665 => x"f8c3c31e",
  2666 => x"c150c048",
  2667 => x"c148dce8",
  2668 => x"c4ffc050",
  2669 => x"c150c048",
  2670 => x"87c9fc49",
  2671 => x"49c0c0c4",
  2672 => x"c287ddfd",
  2673 => x"49bfd4eb",
  2674 => x"c287dcfe",
  2675 => x"49bfd4eb",
  2676 => x"87d6d8fe",
  2677 => x"ecfb49c0",
  2678 => x"49d0c687",
  2679 => x"7087f1f2",
  2680 => x"f7f2494b",
  2681 => x"05987087",
  2682 => x"497387ca",
  2683 => x"7087edf2",
  2684 => x"87f60298",
  2685 => x"ccfb49c1",
  2686 => x"49e4c187",
  2687 => x"7087d1f2",
  2688 => x"d7f2494b",
  2689 => x"05987087",
  2690 => x"497387ca",
  2691 => x"7087cdf2",
  2692 => x"87f60298",
  2693 => x"ecfa49c0",
  2694 => x"2648c087",
  2695 => x"1e4f264b",
  2696 => x"eac21e73",
  2697 => x"c005bffc",
  2698 => x"c9c387ea",
  2699 => x"c4ff49d8",
  2700 => x"b7c087e8",
  2701 => x"87ce04a8",
  2702 => x"49d8c9c3",
  2703 => x"87dac4ff",
  2704 => x"03a8b7c0",
  2705 => x"eac287f2",
  2706 => x"c148bffc",
  2707 => x"c0ebc280",
  2708 => x"87e2c158",
  2709 => x"bffceac2",
  2710 => x"99c1494b",
  2711 => x"87f0c002",
  2712 => x"b7c14973",
  2713 => x"d8ebc229",
  2714 => x"9a4a1181",
  2715 => x"87c6c102",
  2716 => x"06aab7c1",
  2717 => x"1e7287cc",
  2718 => x"49d8c9c3",
  2719 => x"87e6c1ff",
  2720 => x"eac286c4",
  2721 => x"c148bffc",
  2722 => x"c0ebc280",
  2723 => x"87e6c058",
  2724 => x"49d8c9c3",
  2725 => x"87c2c3ff",
  2726 => x"eac24a70",
  2727 => x"87cb02aa",
  2728 => x"02aafac3",
  2729 => x"aac387c5",
  2730 => x"c287cb05",
  2731 => x"48bffcea",
  2732 => x"ebc280c1",
  2733 => x"4b2658c0",
  2734 => x"00004f26",
  2735 => x"00000000",
  2736 => x"00002bf0",
  2737 => x"11141258",
  2738 => x"231c1b1d",
  2739 => x"9194595a",
  2740 => x"f4ebf2f5",
  2741 => x"00002d68",
  2742 => x"f3c8f3ff",
  2743 => x"f250f364",
  2744 => x"1e00f401",
  2745 => x"4b711e73",
  2746 => x"c5e8fe49",
  2747 => x"fcc9c387",
  2748 => x"c702bf97",
  2749 => x"c0c0c487",
  2750 => x"87e4f849",
  2751 => x"e7fe4973",
  2752 => x"4b2687f0",
  2753 => x"731e4f26",
  2754 => x"c34a711e",
  2755 => x"4bbff0c3",
  2756 => x"c5029a72",
  2757 => x"bbc0c287",
  2758 => x"c0c187c3",
  2759 => x"f64973bb",
  2760 => x"f4c787e3",
  2761 => x"87e8ed49",
  2762 => x"ed494b70",
  2763 => x"987087ee",
  2764 => x"7387ca05",
  2765 => x"87e4ed49",
  2766 => x"f6029870",
  2767 => x"264b2687",
  2768 => x"5b5e0e4f",
  2769 => x"4b710e5c",
  2770 => x"d30266cc",
  2771 => x"f0c04c87",
  2772 => x"e9c0028c",
  2773 => x"c1497487",
  2774 => x"e1c00289",
  2775 => x"87f3c087",
  2776 => x"c0029b73",
  2777 => x"c3c387ed",
  2778 => x"c149bff0",
  2779 => x"d4f571b1",
  2780 => x"f7497387",
  2781 => x"497387f1",
  2782 => x"87eed1fe",
  2783 => x"1e7487d5",
  2784 => x"dbf249c0",
  2785 => x"fd497487",
  2786 => x"1e7487fc",
  2787 => x"cff24973",
  2788 => x"c386c887",
  2789 => x"49bff0c3",
  2790 => x"2687eaf4",
  2791 => x"264b264c",
  2792 => x"c4ff1e4f",
  2793 => x"d4ff87df",
  2794 => x"78ffc348",
  2795 => x"87d0dffd",
  2796 => x"cd029870",
  2797 => x"eee8fd87",
  2798 => x"02987087",
  2799 => x"4ac187c4",
  2800 => x"4ac087c2",
  2801 => x"c8029a72",
  2802 => x"ecefc287",
  2803 => x"d6d3fd49",
  2804 => x"fe49c087",
  2805 => x"f787e1f8",
  2806 => x"fbfe87c8",
  2807 => x"fef887e1",
  2808 => x"e5deff87",
  2809 => x"87c1ed87",
  2810 => x"4f2687f4",
  2811 => x"00004b4f",
  2812 => x"72617441",
  2813 => x"54532069",
  2814 => x"30533b3b",
  2815 => x"54532c55",
  2816 => x"6c462c20",
  2817 => x"7970706f",
  2818 => x"3b3a4120",
  2819 => x"2c553153",
  2820 => x"2c205453",
  2821 => x"706f6c46",
  2822 => x"42207970",
  2823 => x"364f3b3a",
  2824 => x"72572c37",
  2825 => x"20657469",
  2826 => x"746f7270",
  2827 => x"2c746365",
  2828 => x"2c66664f",
  2829 => x"422c3a41",
  2830 => x"6f422c3a",
  2831 => x"463b6874",
  2832 => x"474d492c",
  2833 => x"2c4d4f52",
  2834 => x"64616f4c",
  2835 => x"4d4f5220",
  2836 => x"2c31503b",
  2837 => x"43205453",
  2838 => x"69666e6f",
  2839 => x"61727567",
  2840 => x"6e6f6974",
  2841 => x"4f31503b",
  2842 => x"522c3331",
  2843 => x"28204d41",
  2844 => x"6465656e",
  2845 => x"72614820",
  2846 => x"65522064",
  2847 => x"29746573",
  2848 => x"3231352c",
  2849 => x"4d312c4b",
  2850 => x"4d322c42",
  2851 => x"4d342c42",
  2852 => x"4d382c42",
  2853 => x"34312c42",
  2854 => x"503b424d",
  2855 => x"2c384f31",
  2856 => x"65646956",
  2857 => x"6f6d206f",
  2858 => x"4d2c6564",
  2859 => x"2c6f6e6f",
  2860 => x"6f6c6f43",
  2861 => x"503b7275",
  2862 => x"4f4e4f31",
  2863 => x"6968432c",
  2864 => x"74657370",
  2865 => x"2c54532c",
  2866 => x"2c455453",
  2867 => x"6167654d",
  2868 => x"3b455453",
  2869 => x"4a4f3150",
  2870 => x"2054532c",
  2871 => x"74696c42",
  2872 => x"2c726574",
  2873 => x"2c66664f",
  2874 => x"503b6e4f",
  2875 => x"2c4d4f31",
  2876 => x"72657453",
  2877 => x"73206f65",
  2878 => x"646e756f",
  2879 => x"66664f2c",
  2880 => x"3b6e4f2c",
  2881 => x"4b4f3150",
  2882 => x"63532c4c",
  2883 => x"696c6e61",
  2884 => x"2c73656e",
  2885 => x"2c66664f",
  2886 => x"2c253532",
  2887 => x"2c253035",
  2888 => x"3b253537",
  2889 => x"544f3150",
  2890 => x"6d6f432c",
  2891 => x"69736f70",
  2892 => x"62206574",
  2893 => x"646e656c",
  2894 => x"66664f2c",
  2895 => x"3b6e4f2c",
  2896 => x"522c3054",
  2897 => x"74657365",
  2898 => x"6f482820",
  2899 => x"6620646c",
  2900 => x"6820726f",
  2901 => x"20647261",
  2902 => x"65736572",
  2903 => x"563b2974",
  2904 => x"2e33762c",
  2905 => x"002e3034",
  2906 => x"20534f54",
  2907 => x"20202020",
  2908 => x"00474d49",
  2909 => x"00001aaf",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
