
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e8",x"cc",x"c3",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"e8",x"cc",x"c3"),
    18 => (x"48",x"f8",x"f5",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"f8",x"f5",x"c2",x"87"),
    25 => (x"f4",x"f5",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"ec",x"c2",x"87",x"f7"),
    29 => (x"f5",x"c2",x"87",x"eb"),
    30 => (x"f5",x"c2",x"4d",x"f8"),
    31 => (x"ad",x"74",x"4c",x"f8"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"81",x"48",x"73",x"1e"),
    65 => (x"c5",x"02",x"a9",x"73"),
    66 => (x"05",x"53",x"12",x"87"),
    67 => (x"4f",x"26",x"87",x"f6"),
    68 => (x"71",x"1e",x"73",x"1e"),
    69 => (x"4b",x"66",x"c8",x"4a"),
    70 => (x"71",x"8b",x"c1",x"49"),
    71 => (x"87",x"cf",x"02",x"99"),
    72 => (x"d4",x"ff",x"48",x"12"),
    73 => (x"49",x"73",x"78",x"08"),
    74 => (x"99",x"71",x"8b",x"c1"),
    75 => (x"26",x"87",x"f1",x"05"),
    76 => (x"0e",x"4f",x"26",x"4b"),
    77 => (x"0e",x"5c",x"5b",x"5e"),
    78 => (x"d4",x"ff",x"4a",x"71"),
    79 => (x"4b",x"66",x"cc",x"4c"),
    80 => (x"71",x"8b",x"c1",x"49"),
    81 => (x"87",x"ce",x"02",x"99"),
    82 => (x"6c",x"7c",x"ff",x"c3"),
    83 => (x"c1",x"49",x"73",x"52"),
    84 => (x"05",x"99",x"71",x"8b"),
    85 => (x"4c",x"26",x"87",x"f2"),
    86 => (x"4f",x"26",x"4b",x"26"),
    87 => (x"ff",x"1e",x"73",x"1e"),
    88 => (x"ff",x"c3",x"4b",x"d4"),
    89 => (x"c3",x"4a",x"6b",x"7b"),
    90 => (x"49",x"6b",x"7b",x"ff"),
    91 => (x"b1",x"72",x"32",x"c8"),
    92 => (x"6b",x"7b",x"ff",x"c3"),
    93 => (x"71",x"31",x"c8",x"4a"),
    94 => (x"7b",x"ff",x"c3",x"b2"),
    95 => (x"32",x"c8",x"49",x"6b"),
    96 => (x"48",x"71",x"b1",x"72"),
    97 => (x"4f",x"26",x"4b",x"26"),
    98 => (x"5c",x"5b",x"5e",x"0e"),
    99 => (x"4d",x"71",x"0e",x"5d"),
   100 => (x"75",x"4c",x"d4",x"ff"),
   101 => (x"98",x"ff",x"c3",x"48"),
   102 => (x"f5",x"c2",x"7c",x"70"),
   103 => (x"c8",x"05",x"bf",x"f8"),
   104 => (x"48",x"66",x"d0",x"87"),
   105 => (x"a6",x"d4",x"30",x"c9"),
   106 => (x"49",x"66",x"d0",x"58"),
   107 => (x"48",x"71",x"29",x"d8"),
   108 => (x"70",x"98",x"ff",x"c3"),
   109 => (x"49",x"66",x"d0",x"7c"),
   110 => (x"48",x"71",x"29",x"d0"),
   111 => (x"70",x"98",x"ff",x"c3"),
   112 => (x"49",x"66",x"d0",x"7c"),
   113 => (x"48",x"71",x"29",x"c8"),
   114 => (x"70",x"98",x"ff",x"c3"),
   115 => (x"48",x"66",x"d0",x"7c"),
   116 => (x"70",x"98",x"ff",x"c3"),
   117 => (x"d0",x"49",x"75",x"7c"),
   118 => (x"c3",x"48",x"71",x"29"),
   119 => (x"7c",x"70",x"98",x"ff"),
   120 => (x"f0",x"c9",x"4b",x"6c"),
   121 => (x"ff",x"c3",x"4a",x"ff"),
   122 => (x"87",x"cf",x"05",x"ab"),
   123 => (x"6c",x"7c",x"71",x"49"),
   124 => (x"02",x"8a",x"c1",x"4b"),
   125 => (x"ab",x"71",x"87",x"c5"),
   126 => (x"73",x"87",x"f2",x"02"),
   127 => (x"26",x"4d",x"26",x"48"),
   128 => (x"26",x"4b",x"26",x"4c"),
   129 => (x"49",x"c0",x"1e",x"4f"),
   130 => (x"c3",x"48",x"d4",x"ff"),
   131 => (x"81",x"c1",x"78",x"ff"),
   132 => (x"a9",x"b7",x"c8",x"c3"),
   133 => (x"26",x"87",x"f1",x"04"),
   134 => (x"5b",x"5e",x"0e",x"4f"),
   135 => (x"c0",x"0e",x"5d",x"5c"),
   136 => (x"f7",x"c1",x"f0",x"ff"),
   137 => (x"c0",x"c0",x"c1",x"4d"),
   138 => (x"4b",x"c0",x"c0",x"c0"),
   139 => (x"c4",x"87",x"d6",x"ff"),
   140 => (x"c0",x"4c",x"df",x"f8"),
   141 => (x"fd",x"49",x"75",x"1e"),
   142 => (x"86",x"c4",x"87",x"ce"),
   143 => (x"c0",x"05",x"a8",x"c1"),
   144 => (x"d4",x"ff",x"87",x"e5"),
   145 => (x"78",x"ff",x"c3",x"48"),
   146 => (x"e1",x"c0",x"1e",x"73"),
   147 => (x"49",x"e9",x"c1",x"f0"),
   148 => (x"c4",x"87",x"f5",x"fc"),
   149 => (x"05",x"98",x"70",x"86"),
   150 => (x"d4",x"ff",x"87",x"ca"),
   151 => (x"78",x"ff",x"c3",x"48"),
   152 => (x"87",x"cb",x"48",x"c1"),
   153 => (x"c1",x"87",x"de",x"fe"),
   154 => (x"c6",x"ff",x"05",x"8c"),
   155 => (x"26",x"48",x"c0",x"87"),
   156 => (x"26",x"4c",x"26",x"4d"),
   157 => (x"0e",x"4f",x"26",x"4b"),
   158 => (x"0e",x"5c",x"5b",x"5e"),
   159 => (x"c1",x"f0",x"ff",x"c0"),
   160 => (x"d4",x"ff",x"4c",x"c1"),
   161 => (x"78",x"ff",x"c3",x"48"),
   162 => (x"f8",x"49",x"fc",x"ca"),
   163 => (x"4b",x"d3",x"87",x"d9"),
   164 => (x"49",x"74",x"1e",x"c0"),
   165 => (x"c4",x"87",x"f1",x"fb"),
   166 => (x"05",x"98",x"70",x"86"),
   167 => (x"d4",x"ff",x"87",x"ca"),
   168 => (x"78",x"ff",x"c3",x"48"),
   169 => (x"87",x"cb",x"48",x"c1"),
   170 => (x"c1",x"87",x"da",x"fd"),
   171 => (x"df",x"ff",x"05",x"8b"),
   172 => (x"26",x"48",x"c0",x"87"),
   173 => (x"26",x"4b",x"26",x"4c"),
   174 => (x"00",x"00",x"00",x"4f"),
   175 => (x"00",x"44",x"4d",x"43"),
   176 => (x"43",x"48",x"44",x"53"),
   177 => (x"69",x"61",x"66",x"20"),
   178 => (x"00",x"0a",x"21",x"6c"),
   179 => (x"52",x"52",x"45",x"49"),
   180 => (x"00",x"00",x"00",x"00"),
   181 => (x"00",x"49",x"50",x"53"),
   182 => (x"74",x"69",x"72",x"57"),
   183 => (x"61",x"66",x"20",x"65"),
   184 => (x"64",x"65",x"6c",x"69"),
   185 => (x"5e",x"0e",x"00",x"0a"),
   186 => (x"0e",x"5d",x"5c",x"5b"),
   187 => (x"ff",x"4d",x"ff",x"c3"),
   188 => (x"d0",x"fc",x"4b",x"d4"),
   189 => (x"1e",x"ea",x"c6",x"87"),
   190 => (x"c1",x"f0",x"e1",x"c0"),
   191 => (x"c7",x"fa",x"49",x"c8"),
   192 => (x"c1",x"86",x"c4",x"87"),
   193 => (x"87",x"c8",x"02",x"a8"),
   194 => (x"c0",x"87",x"ec",x"fd"),
   195 => (x"87",x"e8",x"c1",x"48"),
   196 => (x"70",x"87",x"c9",x"f9"),
   197 => (x"ff",x"ff",x"cf",x"49"),
   198 => (x"a9",x"ea",x"c6",x"99"),
   199 => (x"fd",x"87",x"c8",x"02"),
   200 => (x"48",x"c0",x"87",x"d5"),
   201 => (x"75",x"87",x"d1",x"c1"),
   202 => (x"4c",x"f1",x"c0",x"7b"),
   203 => (x"70",x"87",x"ea",x"fb"),
   204 => (x"ec",x"c0",x"02",x"98"),
   205 => (x"c0",x"1e",x"c0",x"87"),
   206 => (x"fa",x"c1",x"f0",x"ff"),
   207 => (x"87",x"c8",x"f9",x"49"),
   208 => (x"98",x"70",x"86",x"c4"),
   209 => (x"75",x"87",x"da",x"05"),
   210 => (x"75",x"49",x"6b",x"7b"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"c1",x"7b",x"75",x"7b"),
   213 => (x"c4",x"02",x"99",x"c0"),
   214 => (x"db",x"48",x"c1",x"87"),
   215 => (x"d7",x"48",x"c0",x"87"),
   216 => (x"05",x"ac",x"c2",x"87"),
   217 => (x"c0",x"cb",x"87",x"ca"),
   218 => (x"87",x"fb",x"f4",x"49"),
   219 => (x"87",x"c8",x"48",x"c0"),
   220 => (x"fe",x"05",x"8c",x"c1"),
   221 => (x"48",x"c0",x"87",x"f6"),
   222 => (x"4c",x"26",x"4d",x"26"),
   223 => (x"4f",x"26",x"4b",x"26"),
   224 => (x"5c",x"5b",x"5e",x"0e"),
   225 => (x"d0",x"ff",x"0e",x"5d"),
   226 => (x"d0",x"e5",x"c0",x"4d"),
   227 => (x"c2",x"4c",x"c0",x"c1"),
   228 => (x"c1",x"48",x"f8",x"f5"),
   229 => (x"49",x"d4",x"cb",x"78"),
   230 => (x"c7",x"87",x"cc",x"f4"),
   231 => (x"f9",x"7d",x"c2",x"4b"),
   232 => (x"7d",x"c3",x"87",x"e3"),
   233 => (x"49",x"74",x"1e",x"c0"),
   234 => (x"c4",x"87",x"dd",x"f7"),
   235 => (x"05",x"a8",x"c1",x"86"),
   236 => (x"c2",x"4b",x"87",x"c1"),
   237 => (x"87",x"cb",x"05",x"ab"),
   238 => (x"f3",x"49",x"cc",x"cb"),
   239 => (x"48",x"c0",x"87",x"e9"),
   240 => (x"c1",x"87",x"f6",x"c0"),
   241 => (x"d4",x"ff",x"05",x"8b"),
   242 => (x"87",x"da",x"fc",x"87"),
   243 => (x"58",x"fc",x"f5",x"c2"),
   244 => (x"cd",x"05",x"98",x"70"),
   245 => (x"c0",x"1e",x"c1",x"87"),
   246 => (x"d0",x"c1",x"f0",x"ff"),
   247 => (x"87",x"e8",x"f6",x"49"),
   248 => (x"d4",x"ff",x"86",x"c4"),
   249 => (x"78",x"ff",x"c3",x"48"),
   250 => (x"c2",x"87",x"ee",x"c4"),
   251 => (x"c2",x"58",x"c0",x"f6"),
   252 => (x"48",x"d4",x"ff",x"7d"),
   253 => (x"c1",x"78",x"ff",x"c3"),
   254 => (x"26",x"4d",x"26",x"48"),
   255 => (x"26",x"4b",x"26",x"4c"),
   256 => (x"5b",x"5e",x"0e",x"4f"),
   257 => (x"71",x"0e",x"5d",x"5c"),
   258 => (x"4c",x"ff",x"c3",x"4d"),
   259 => (x"74",x"4b",x"d4",x"ff"),
   260 => (x"48",x"d0",x"ff",x"7b"),
   261 => (x"74",x"78",x"c3",x"c4"),
   262 => (x"c0",x"1e",x"75",x"7b"),
   263 => (x"d8",x"c1",x"f0",x"ff"),
   264 => (x"87",x"e4",x"f5",x"49"),
   265 => (x"98",x"70",x"86",x"c4"),
   266 => (x"cb",x"87",x"cb",x"02"),
   267 => (x"f6",x"f1",x"49",x"d8"),
   268 => (x"c0",x"48",x"c1",x"87"),
   269 => (x"7b",x"74",x"87",x"ee"),
   270 => (x"c8",x"7b",x"fe",x"c3"),
   271 => (x"66",x"d4",x"1e",x"c0"),
   272 => (x"87",x"cc",x"f3",x"49"),
   273 => (x"7b",x"74",x"86",x"c4"),
   274 => (x"7b",x"74",x"7b",x"74"),
   275 => (x"4a",x"e0",x"da",x"d8"),
   276 => (x"05",x"6b",x"7b",x"74"),
   277 => (x"8a",x"c1",x"87",x"c5"),
   278 => (x"74",x"87",x"f5",x"05"),
   279 => (x"48",x"d0",x"ff",x"7b"),
   280 => (x"48",x"c0",x"78",x"c2"),
   281 => (x"4c",x"26",x"4d",x"26"),
   282 => (x"4f",x"26",x"4b",x"26"),
   283 => (x"5c",x"5b",x"5e",x"0e"),
   284 => (x"86",x"fc",x"0e",x"5d"),
   285 => (x"d4",x"ff",x"4b",x"71"),
   286 => (x"c5",x"7e",x"c0",x"4c"),
   287 => (x"4a",x"df",x"cd",x"ee"),
   288 => (x"6c",x"7c",x"ff",x"c3"),
   289 => (x"a8",x"fe",x"c3",x"48"),
   290 => (x"87",x"f8",x"c0",x"05"),
   291 => (x"9b",x"73",x"4d",x"74"),
   292 => (x"d4",x"87",x"cc",x"02"),
   293 => (x"49",x"73",x"1e",x"66"),
   294 => (x"c4",x"87",x"d8",x"f2"),
   295 => (x"ff",x"87",x"d4",x"86"),
   296 => (x"d1",x"c4",x"48",x"d0"),
   297 => (x"4a",x"66",x"d4",x"78"),
   298 => (x"c1",x"7d",x"ff",x"c3"),
   299 => (x"87",x"f8",x"05",x"8a"),
   300 => (x"c3",x"5a",x"a6",x"d8"),
   301 => (x"73",x"7c",x"7c",x"ff"),
   302 => (x"87",x"c5",x"05",x"9b"),
   303 => (x"d0",x"48",x"d0",x"ff"),
   304 => (x"7e",x"4a",x"c1",x"78"),
   305 => (x"fe",x"05",x"8a",x"c1"),
   306 => (x"48",x"6e",x"87",x"f6"),
   307 => (x"4d",x"26",x"8e",x"fc"),
   308 => (x"4b",x"26",x"4c",x"26"),
   309 => (x"73",x"1e",x"4f",x"26"),
   310 => (x"c0",x"4a",x"71",x"1e"),
   311 => (x"48",x"d4",x"ff",x"4b"),
   312 => (x"ff",x"78",x"ff",x"c3"),
   313 => (x"c3",x"c4",x"48",x"d0"),
   314 => (x"48",x"d4",x"ff",x"78"),
   315 => (x"72",x"78",x"ff",x"c3"),
   316 => (x"f0",x"ff",x"c0",x"1e"),
   317 => (x"f2",x"49",x"d1",x"c1"),
   318 => (x"86",x"c4",x"87",x"ce"),
   319 => (x"d2",x"05",x"98",x"70"),
   320 => (x"1e",x"c0",x"c8",x"87"),
   321 => (x"fd",x"49",x"66",x"cc"),
   322 => (x"86",x"c4",x"87",x"e2"),
   323 => (x"d0",x"ff",x"4b",x"70"),
   324 => (x"73",x"78",x"c2",x"48"),
   325 => (x"26",x"4b",x"26",x"48"),
   326 => (x"5b",x"5e",x"0e",x"4f"),
   327 => (x"c0",x"0e",x"5d",x"5c"),
   328 => (x"f0",x"ff",x"c0",x"1e"),
   329 => (x"f1",x"49",x"c9",x"c1"),
   330 => (x"1e",x"d2",x"87",x"de"),
   331 => (x"49",x"c8",x"f6",x"c2"),
   332 => (x"c8",x"87",x"f9",x"fc"),
   333 => (x"c1",x"4c",x"c0",x"86"),
   334 => (x"ac",x"b7",x"d2",x"84"),
   335 => (x"c2",x"87",x"f8",x"04"),
   336 => (x"bf",x"97",x"c8",x"f6"),
   337 => (x"99",x"c0",x"c3",x"49"),
   338 => (x"05",x"a9",x"c0",x"c1"),
   339 => (x"c2",x"87",x"e7",x"c0"),
   340 => (x"bf",x"97",x"cf",x"f6"),
   341 => (x"c2",x"31",x"d0",x"49"),
   342 => (x"bf",x"97",x"d0",x"f6"),
   343 => (x"72",x"32",x"c8",x"4a"),
   344 => (x"d1",x"f6",x"c2",x"b1"),
   345 => (x"b1",x"4a",x"bf",x"97"),
   346 => (x"ff",x"cf",x"4c",x"71"),
   347 => (x"c1",x"9c",x"ff",x"ff"),
   348 => (x"c1",x"34",x"ca",x"84"),
   349 => (x"f6",x"c2",x"87",x"e7"),
   350 => (x"49",x"bf",x"97",x"d1"),
   351 => (x"99",x"c6",x"31",x"c1"),
   352 => (x"97",x"d2",x"f6",x"c2"),
   353 => (x"b7",x"c7",x"4a",x"bf"),
   354 => (x"c2",x"b1",x"72",x"2a"),
   355 => (x"bf",x"97",x"cd",x"f6"),
   356 => (x"9d",x"cf",x"4d",x"4a"),
   357 => (x"97",x"ce",x"f6",x"c2"),
   358 => (x"9a",x"c3",x"4a",x"bf"),
   359 => (x"f6",x"c2",x"32",x"ca"),
   360 => (x"4b",x"bf",x"97",x"cf"),
   361 => (x"b2",x"73",x"33",x"c2"),
   362 => (x"97",x"d0",x"f6",x"c2"),
   363 => (x"c0",x"c3",x"4b",x"bf"),
   364 => (x"2b",x"b7",x"c6",x"9b"),
   365 => (x"81",x"c2",x"b2",x"73"),
   366 => (x"30",x"71",x"48",x"c1"),
   367 => (x"48",x"c1",x"49",x"70"),
   368 => (x"4d",x"70",x"30",x"75"),
   369 => (x"84",x"c1",x"4c",x"72"),
   370 => (x"c0",x"c8",x"94",x"71"),
   371 => (x"cc",x"06",x"ad",x"b7"),
   372 => (x"b7",x"34",x"c1",x"87"),
   373 => (x"b7",x"c0",x"c8",x"2d"),
   374 => (x"f4",x"ff",x"01",x"ad"),
   375 => (x"26",x"48",x"74",x"87"),
   376 => (x"26",x"4c",x"26",x"4d"),
   377 => (x"0e",x"4f",x"26",x"4b"),
   378 => (x"5d",x"5c",x"5b",x"5e"),
   379 => (x"c2",x"86",x"fc",x"0e"),
   380 => (x"c0",x"48",x"f0",x"fe"),
   381 => (x"e8",x"f6",x"c2",x"78"),
   382 => (x"fb",x"49",x"c0",x"1e"),
   383 => (x"86",x"c4",x"87",x"d8"),
   384 => (x"c5",x"05",x"98",x"70"),
   385 => (x"c9",x"48",x"c0",x"87"),
   386 => (x"4d",x"c0",x"87",x"d2"),
   387 => (x"48",x"ec",x"c3",x"c3"),
   388 => (x"f7",x"c2",x"78",x"c1"),
   389 => (x"e1",x"c0",x"4a",x"de"),
   390 => (x"4b",x"c8",x"49",x"f4"),
   391 => (x"70",x"87",x"c7",x"eb"),
   392 => (x"87",x"c6",x"05",x"98"),
   393 => (x"48",x"ec",x"c3",x"c3"),
   394 => (x"f7",x"c2",x"78",x"c0"),
   395 => (x"e2",x"c0",x"4a",x"fa"),
   396 => (x"4b",x"c8",x"49",x"c0"),
   397 => (x"70",x"87",x"ef",x"ea"),
   398 => (x"87",x"c6",x"05",x"98"),
   399 => (x"48",x"ec",x"c3",x"c3"),
   400 => (x"c3",x"c3",x"78",x"c0"),
   401 => (x"c0",x"02",x"bf",x"ec"),
   402 => (x"fd",x"c2",x"87",x"fd"),
   403 => (x"c2",x"4d",x"bf",x"ee"),
   404 => (x"bf",x"9f",x"e6",x"fe"),
   405 => (x"d6",x"c5",x"48",x"7e"),
   406 => (x"c7",x"05",x"a8",x"ea"),
   407 => (x"ee",x"fd",x"c2",x"87"),
   408 => (x"87",x"ce",x"4d",x"bf"),
   409 => (x"e9",x"ca",x"48",x"6e"),
   410 => (x"c5",x"02",x"a8",x"d5"),
   411 => (x"c7",x"48",x"c0",x"87"),
   412 => (x"f6",x"c2",x"87",x"ea"),
   413 => (x"49",x"75",x"1e",x"e8"),
   414 => (x"c4",x"87",x"db",x"f9"),
   415 => (x"05",x"98",x"70",x"86"),
   416 => (x"48",x"c0",x"87",x"c5"),
   417 => (x"c2",x"87",x"d5",x"c7"),
   418 => (x"c0",x"4a",x"fa",x"f7"),
   419 => (x"c8",x"49",x"cc",x"e2"),
   420 => (x"87",x"d2",x"e9",x"4b"),
   421 => (x"c8",x"05",x"98",x"70"),
   422 => (x"f0",x"fe",x"c2",x"87"),
   423 => (x"d8",x"78",x"c1",x"48"),
   424 => (x"de",x"f7",x"c2",x"87"),
   425 => (x"d8",x"e2",x"c0",x"4a"),
   426 => (x"e8",x"4b",x"c8",x"49"),
   427 => (x"98",x"70",x"87",x"f8"),
   428 => (x"87",x"c5",x"c0",x"02"),
   429 => (x"e3",x"c6",x"48",x"c0"),
   430 => (x"e6",x"fe",x"c2",x"87"),
   431 => (x"c1",x"49",x"bf",x"97"),
   432 => (x"c0",x"05",x"a9",x"d5"),
   433 => (x"fe",x"c2",x"87",x"cd"),
   434 => (x"49",x"bf",x"97",x"e7"),
   435 => (x"02",x"a9",x"ea",x"c2"),
   436 => (x"c0",x"87",x"c5",x"c0"),
   437 => (x"87",x"c4",x"c6",x"48"),
   438 => (x"97",x"e8",x"f6",x"c2"),
   439 => (x"c3",x"48",x"7e",x"bf"),
   440 => (x"c0",x"02",x"a8",x"e9"),
   441 => (x"48",x"6e",x"87",x"ce"),
   442 => (x"02",x"a8",x"eb",x"c3"),
   443 => (x"c0",x"87",x"c5",x"c0"),
   444 => (x"87",x"e8",x"c5",x"48"),
   445 => (x"97",x"f3",x"f6",x"c2"),
   446 => (x"05",x"99",x"49",x"bf"),
   447 => (x"c2",x"87",x"cc",x"c0"),
   448 => (x"bf",x"97",x"f4",x"f6"),
   449 => (x"02",x"a9",x"c2",x"49"),
   450 => (x"c0",x"87",x"c5",x"c0"),
   451 => (x"87",x"cc",x"c5",x"48"),
   452 => (x"97",x"f5",x"f6",x"c2"),
   453 => (x"fe",x"c2",x"48",x"bf"),
   454 => (x"4c",x"70",x"58",x"ec"),
   455 => (x"c2",x"88",x"c1",x"48"),
   456 => (x"c2",x"58",x"f0",x"fe"),
   457 => (x"bf",x"97",x"f6",x"f6"),
   458 => (x"c2",x"81",x"75",x"49"),
   459 => (x"bf",x"97",x"f7",x"f6"),
   460 => (x"72",x"32",x"c8",x"4a"),
   461 => (x"c3",x"c3",x"7e",x"a1"),
   462 => (x"78",x"6e",x"48",x"c8"),
   463 => (x"97",x"f8",x"f6",x"c2"),
   464 => (x"c3",x"c3",x"48",x"bf"),
   465 => (x"fe",x"c2",x"58",x"e0"),
   466 => (x"c2",x"02",x"bf",x"f0"),
   467 => (x"f7",x"c2",x"87",x"d3"),
   468 => (x"e1",x"c0",x"4a",x"fa"),
   469 => (x"4b",x"c8",x"49",x"e8"),
   470 => (x"70",x"87",x"cb",x"e6"),
   471 => (x"c5",x"c0",x"02",x"98"),
   472 => (x"c3",x"48",x"c0",x"87"),
   473 => (x"fe",x"c2",x"87",x"f6"),
   474 => (x"c3",x"4c",x"bf",x"e8"),
   475 => (x"c2",x"5c",x"dc",x"c3"),
   476 => (x"bf",x"97",x"cd",x"f7"),
   477 => (x"c2",x"31",x"c8",x"49"),
   478 => (x"bf",x"97",x"cc",x"f7"),
   479 => (x"c2",x"49",x"a1",x"4a"),
   480 => (x"bf",x"97",x"ce",x"f7"),
   481 => (x"72",x"32",x"d0",x"4a"),
   482 => (x"f7",x"c2",x"49",x"a1"),
   483 => (x"4a",x"bf",x"97",x"cf"),
   484 => (x"a1",x"72",x"32",x"d8"),
   485 => (x"e4",x"c3",x"c3",x"49"),
   486 => (x"dc",x"c3",x"c3",x"59"),
   487 => (x"c3",x"c3",x"91",x"bf"),
   488 => (x"c3",x"81",x"bf",x"c8"),
   489 => (x"c2",x"59",x"d0",x"c3"),
   490 => (x"bf",x"97",x"d5",x"f7"),
   491 => (x"c2",x"32",x"c8",x"4a"),
   492 => (x"bf",x"97",x"d4",x"f7"),
   493 => (x"c2",x"4a",x"a2",x"4b"),
   494 => (x"bf",x"97",x"d6",x"f7"),
   495 => (x"73",x"33",x"d0",x"4b"),
   496 => (x"f7",x"c2",x"4a",x"a2"),
   497 => (x"4b",x"bf",x"97",x"d7"),
   498 => (x"33",x"d8",x"9b",x"cf"),
   499 => (x"c3",x"4a",x"a2",x"73"),
   500 => (x"c2",x"5a",x"d4",x"c3"),
   501 => (x"c3",x"92",x"74",x"8a"),
   502 => (x"72",x"48",x"d4",x"c3"),
   503 => (x"c7",x"c1",x"78",x"a1"),
   504 => (x"fa",x"f6",x"c2",x"87"),
   505 => (x"c8",x"49",x"bf",x"97"),
   506 => (x"f9",x"f6",x"c2",x"31"),
   507 => (x"a1",x"4a",x"bf",x"97"),
   508 => (x"c7",x"31",x"c5",x"49"),
   509 => (x"29",x"c9",x"81",x"ff"),
   510 => (x"59",x"dc",x"c3",x"c3"),
   511 => (x"97",x"ff",x"f6",x"c2"),
   512 => (x"32",x"c8",x"4a",x"bf"),
   513 => (x"97",x"fe",x"f6",x"c2"),
   514 => (x"4a",x"a2",x"4b",x"bf"),
   515 => (x"5a",x"e4",x"c3",x"c3"),
   516 => (x"bf",x"dc",x"c3",x"c3"),
   517 => (x"c3",x"82",x"6e",x"92"),
   518 => (x"c3",x"5a",x"d8",x"c3"),
   519 => (x"c0",x"48",x"d0",x"c3"),
   520 => (x"cc",x"c3",x"c3",x"78"),
   521 => (x"78",x"a1",x"72",x"48"),
   522 => (x"48",x"e4",x"c3",x"c3"),
   523 => (x"bf",x"d0",x"c3",x"c3"),
   524 => (x"e8",x"c3",x"c3",x"78"),
   525 => (x"d4",x"c3",x"c3",x"48"),
   526 => (x"fe",x"c2",x"78",x"bf"),
   527 => (x"c0",x"02",x"bf",x"f0"),
   528 => (x"48",x"74",x"87",x"c9"),
   529 => (x"7e",x"70",x"30",x"c4"),
   530 => (x"c3",x"87",x"c9",x"c0"),
   531 => (x"48",x"bf",x"d8",x"c3"),
   532 => (x"7e",x"70",x"30",x"c4"),
   533 => (x"48",x"f4",x"fe",x"c2"),
   534 => (x"48",x"c1",x"78",x"6e"),
   535 => (x"4d",x"26",x"8e",x"fc"),
   536 => (x"4b",x"26",x"4c",x"26"),
   537 => (x"00",x"00",x"4f",x"26"),
   538 => (x"33",x"54",x"41",x"46"),
   539 => (x"20",x"20",x"20",x"32"),
   540 => (x"00",x"00",x"00",x"00"),
   541 => (x"31",x"54",x"41",x"46"),
   542 => (x"20",x"20",x"20",x"36"),
   543 => (x"00",x"00",x"00",x"00"),
   544 => (x"33",x"54",x"41",x"46"),
   545 => (x"20",x"20",x"20",x"32"),
   546 => (x"00",x"00",x"00",x"00"),
   547 => (x"33",x"54",x"41",x"46"),
   548 => (x"20",x"20",x"20",x"32"),
   549 => (x"00",x"00",x"00",x"00"),
   550 => (x"31",x"54",x"41",x"46"),
   551 => (x"20",x"20",x"20",x"36"),
   552 => (x"5b",x"5e",x"0e",x"00"),
   553 => (x"71",x"0e",x"5d",x"5c"),
   554 => (x"f0",x"fe",x"c2",x"4a"),
   555 => (x"87",x"cb",x"02",x"bf"),
   556 => (x"2b",x"c7",x"4b",x"72"),
   557 => (x"ff",x"c1",x"4d",x"72"),
   558 => (x"72",x"87",x"c9",x"9d"),
   559 => (x"72",x"2b",x"c8",x"4b"),
   560 => (x"9d",x"ff",x"c3",x"4d"),
   561 => (x"bf",x"c8",x"c3",x"c3"),
   562 => (x"e8",x"f9",x"c0",x"83"),
   563 => (x"d9",x"02",x"ab",x"bf"),
   564 => (x"ec",x"f9",x"c0",x"87"),
   565 => (x"e8",x"f6",x"c2",x"5b"),
   566 => (x"ef",x"49",x"73",x"1e"),
   567 => (x"86",x"c4",x"87",x"f8"),
   568 => (x"c5",x"05",x"98",x"70"),
   569 => (x"c0",x"48",x"c0",x"87"),
   570 => (x"fe",x"c2",x"87",x"e6"),
   571 => (x"d2",x"02",x"bf",x"f0"),
   572 => (x"c4",x"49",x"75",x"87"),
   573 => (x"e8",x"f6",x"c2",x"91"),
   574 => (x"cf",x"4c",x"69",x"81"),
   575 => (x"ff",x"ff",x"ff",x"ff"),
   576 => (x"75",x"87",x"cb",x"9c"),
   577 => (x"c2",x"91",x"c2",x"49"),
   578 => (x"9f",x"81",x"e8",x"f6"),
   579 => (x"48",x"74",x"4c",x"69"),
   580 => (x"4c",x"26",x"4d",x"26"),
   581 => (x"4f",x"26",x"4b",x"26"),
   582 => (x"5c",x"5b",x"5e",x"0e"),
   583 => (x"86",x"f4",x"0e",x"5d"),
   584 => (x"c4",x"59",x"a6",x"c8"),
   585 => (x"80",x"c8",x"48",x"66"),
   586 => (x"c0",x"48",x"7e",x"70"),
   587 => (x"49",x"c1",x"1e",x"78"),
   588 => (x"87",x"f9",x"cc",x"49"),
   589 => (x"4c",x"70",x"86",x"c4"),
   590 => (x"fc",x"c0",x"02",x"9c"),
   591 => (x"f8",x"fe",x"c2",x"87"),
   592 => (x"49",x"66",x"dc",x"4a"),
   593 => (x"87",x"c3",x"de",x"ff"),
   594 => (x"c0",x"02",x"98",x"70"),
   595 => (x"4a",x"74",x"87",x"eb"),
   596 => (x"cb",x"49",x"66",x"dc"),
   597 => (x"cd",x"de",x"ff",x"4b"),
   598 => (x"02",x"98",x"70",x"87"),
   599 => (x"1e",x"c0",x"87",x"db"),
   600 => (x"c4",x"02",x"9c",x"74"),
   601 => (x"c2",x"4d",x"c0",x"87"),
   602 => (x"75",x"4d",x"c1",x"87"),
   603 => (x"87",x"fd",x"cb",x"49"),
   604 => (x"4c",x"70",x"86",x"c4"),
   605 => (x"c4",x"ff",x"05",x"9c"),
   606 => (x"02",x"9c",x"74",x"87"),
   607 => (x"dc",x"87",x"f4",x"c1"),
   608 => (x"48",x"6e",x"49",x"a4"),
   609 => (x"a4",x"da",x"78",x"69"),
   610 => (x"4d",x"66",x"c4",x"49"),
   611 => (x"69",x"9f",x"85",x"c4"),
   612 => (x"f0",x"fe",x"c2",x"7d"),
   613 => (x"87",x"d2",x"02",x"bf"),
   614 => (x"9f",x"49",x"a4",x"d4"),
   615 => (x"ff",x"c0",x"49",x"69"),
   616 => (x"48",x"71",x"99",x"ff"),
   617 => (x"7e",x"70",x"30",x"d0"),
   618 => (x"7e",x"c0",x"87",x"c2"),
   619 => (x"6d",x"48",x"49",x"6e"),
   620 => (x"c4",x"7d",x"70",x"80"),
   621 => (x"78",x"c0",x"48",x"66"),
   622 => (x"cc",x"49",x"66",x"c4"),
   623 => (x"c4",x"79",x"6d",x"81"),
   624 => (x"81",x"d0",x"49",x"66"),
   625 => (x"a6",x"c8",x"79",x"c0"),
   626 => (x"c8",x"78",x"c0",x"48"),
   627 => (x"66",x"c4",x"4c",x"66"),
   628 => (x"74",x"82",x"d4",x"4a"),
   629 => (x"72",x"91",x"c8",x"49"),
   630 => (x"41",x"c0",x"49",x"a1"),
   631 => (x"84",x"c1",x"79",x"6d"),
   632 => (x"04",x"ac",x"b7",x"c6"),
   633 => (x"c4",x"87",x"e7",x"ff"),
   634 => (x"c4",x"c1",x"49",x"66"),
   635 => (x"c1",x"79",x"c0",x"81"),
   636 => (x"c0",x"87",x"c2",x"48"),
   637 => (x"26",x"8e",x"f4",x"48"),
   638 => (x"26",x"4c",x"26",x"4d"),
   639 => (x"0e",x"4f",x"26",x"4b"),
   640 => (x"5d",x"5c",x"5b",x"5e"),
   641 => (x"d0",x"4c",x"71",x"0e"),
   642 => (x"6c",x"4a",x"4d",x"66"),
   643 => (x"4d",x"a1",x"72",x"49"),
   644 => (x"ec",x"fe",x"c2",x"b9"),
   645 => (x"ba",x"ff",x"4a",x"bf"),
   646 => (x"99",x"71",x"99",x"72"),
   647 => (x"87",x"e4",x"c0",x"02"),
   648 => (x"6b",x"4b",x"a4",x"c4"),
   649 => (x"87",x"f9",x"f9",x"49"),
   650 => (x"fe",x"c2",x"7b",x"70"),
   651 => (x"6c",x"49",x"bf",x"e8"),
   652 => (x"75",x"7c",x"71",x"81"),
   653 => (x"ec",x"fe",x"c2",x"b9"),
   654 => (x"ba",x"ff",x"4a",x"bf"),
   655 => (x"99",x"71",x"99",x"72"),
   656 => (x"87",x"dc",x"ff",x"05"),
   657 => (x"4d",x"26",x"7c",x"75"),
   658 => (x"4b",x"26",x"4c",x"26"),
   659 => (x"73",x"1e",x"4f",x"26"),
   660 => (x"c3",x"4b",x"71",x"1e"),
   661 => (x"49",x"bf",x"cc",x"c3"),
   662 => (x"6a",x"4a",x"a3",x"c4"),
   663 => (x"c2",x"8a",x"c2",x"4a"),
   664 => (x"92",x"bf",x"e8",x"fe"),
   665 => (x"c2",x"49",x"a1",x"72"),
   666 => (x"4a",x"bf",x"ec",x"fe"),
   667 => (x"a1",x"72",x"9a",x"6b"),
   668 => (x"ec",x"f9",x"c0",x"49"),
   669 => (x"1e",x"66",x"c8",x"59"),
   670 => (x"87",x"da",x"e9",x"71"),
   671 => (x"98",x"70",x"86",x"c4"),
   672 => (x"c0",x"87",x"c4",x"05"),
   673 => (x"c1",x"87",x"c2",x"48"),
   674 => (x"26",x"4b",x"26",x"48"),
   675 => (x"1e",x"73",x"1e",x"4f"),
   676 => (x"c3",x"c3",x"4b",x"71"),
   677 => (x"c4",x"49",x"bf",x"cc"),
   678 => (x"4a",x"6a",x"4a",x"a3"),
   679 => (x"fe",x"c2",x"8a",x"c2"),
   680 => (x"72",x"92",x"bf",x"e8"),
   681 => (x"fe",x"c2",x"49",x"a1"),
   682 => (x"6b",x"4a",x"bf",x"ec"),
   683 => (x"49",x"a1",x"72",x"9a"),
   684 => (x"59",x"ec",x"f9",x"c0"),
   685 => (x"71",x"1e",x"66",x"c8"),
   686 => (x"c4",x"87",x"c6",x"e5"),
   687 => (x"05",x"98",x"70",x"86"),
   688 => (x"48",x"c0",x"87",x"c4"),
   689 => (x"48",x"c1",x"87",x"c2"),
   690 => (x"4f",x"26",x"4b",x"26"),
   691 => (x"5c",x"5b",x"5e",x"0e"),
   692 => (x"86",x"e0",x"0e",x"5d"),
   693 => (x"f0",x"c0",x"4b",x"71"),
   694 => (x"29",x"c9",x"49",x"66"),
   695 => (x"c2",x"59",x"a6",x"c8"),
   696 => (x"49",x"bf",x"ec",x"fe"),
   697 => (x"4a",x"71",x"b9",x"ff"),
   698 => (x"d8",x"9a",x"66",x"c4"),
   699 => (x"99",x"6b",x"5a",x"a6"),
   700 => (x"c4",x"59",x"a6",x"d0"),
   701 => (x"a6",x"d0",x"7e",x"a3"),
   702 => (x"78",x"bf",x"6e",x"48"),
   703 => (x"cc",x"48",x"66",x"d4"),
   704 => (x"c6",x"05",x"a8",x"66"),
   705 => (x"7b",x"66",x"c4",x"87"),
   706 => (x"d8",x"87",x"c1",x"c3"),
   707 => (x"ff",x"c1",x"48",x"a6"),
   708 => (x"ff",x"ff",x"ff",x"ff"),
   709 => (x"ff",x"80",x"c4",x"78"),
   710 => (x"c8",x"4c",x"c0",x"78"),
   711 => (x"a3",x"d4",x"48",x"a6"),
   712 => (x"c8",x"49",x"74",x"78"),
   713 => (x"81",x"66",x"c8",x"91"),
   714 => (x"4d",x"4a",x"66",x"d4"),
   715 => (x"b7",x"c0",x"8d",x"69"),
   716 => (x"87",x"ce",x"04",x"ad"),
   717 => (x"ad",x"b7",x"66",x"d8"),
   718 => (x"c0",x"87",x"c7",x"03"),
   719 => (x"dc",x"5c",x"a6",x"e0"),
   720 => (x"84",x"c1",x"5d",x"a6"),
   721 => (x"04",x"ac",x"b7",x"c6"),
   722 => (x"dc",x"87",x"d0",x"ff"),
   723 => (x"b7",x"c0",x"48",x"66"),
   724 => (x"87",x"d0",x"04",x"a8"),
   725 => (x"c8",x"49",x"66",x"dc"),
   726 => (x"81",x"66",x"c8",x"91"),
   727 => (x"48",x"6e",x"7b",x"21"),
   728 => (x"87",x"c9",x"78",x"69"),
   729 => (x"a3",x"cc",x"7b",x"c0"),
   730 => (x"69",x"48",x"6e",x"49"),
   731 => (x"48",x"66",x"c4",x"78"),
   732 => (x"a6",x"c8",x"88",x"6b"),
   733 => (x"e8",x"fe",x"c2",x"58"),
   734 => (x"90",x"c8",x"48",x"bf"),
   735 => (x"66",x"c4",x"7e",x"70"),
   736 => (x"01",x"a8",x"6e",x"48"),
   737 => (x"66",x"c4",x"87",x"c9"),
   738 => (x"03",x"a8",x"6e",x"48"),
   739 => (x"c1",x"87",x"f3",x"c0"),
   740 => (x"6a",x"4a",x"a3",x"c4"),
   741 => (x"c8",x"91",x"c8",x"49"),
   742 => (x"66",x"cc",x"81",x"66"),
   743 => (x"c8",x"49",x"6a",x"79"),
   744 => (x"81",x"66",x"c8",x"91"),
   745 => (x"66",x"d0",x"81",x"c4"),
   746 => (x"48",x"7e",x"6a",x"79"),
   747 => (x"c7",x"05",x"a8",x"c5"),
   748 => (x"48",x"a6",x"c8",x"87"),
   749 => (x"87",x"c7",x"78",x"c0"),
   750 => (x"80",x"c1",x"48",x"6e"),
   751 => (x"c8",x"58",x"a6",x"cc"),
   752 => (x"66",x"c4",x"7a",x"66"),
   753 => (x"f8",x"49",x"73",x"1e"),
   754 => (x"86",x"c4",x"87",x"f5"),
   755 => (x"1e",x"e8",x"f6",x"c2"),
   756 => (x"f9",x"f9",x"49",x"73"),
   757 => (x"49",x"a3",x"d0",x"87"),
   758 => (x"79",x"66",x"f4",x"c0"),
   759 => (x"26",x"8e",x"dc",x"ff"),
   760 => (x"26",x"4c",x"26",x"4d"),
   761 => (x"0e",x"4f",x"26",x"4b"),
   762 => (x"0e",x"5c",x"5b",x"5e"),
   763 => (x"4b",x"c0",x"4a",x"71"),
   764 => (x"c0",x"02",x"9a",x"72"),
   765 => (x"a2",x"da",x"87",x"e0"),
   766 => (x"4b",x"69",x"9f",x"49"),
   767 => (x"bf",x"f0",x"fe",x"c2"),
   768 => (x"d4",x"87",x"cf",x"02"),
   769 => (x"69",x"9f",x"49",x"a2"),
   770 => (x"ff",x"c0",x"4c",x"49"),
   771 => (x"34",x"d0",x"9c",x"ff"),
   772 => (x"4c",x"c0",x"87",x"c2"),
   773 => (x"9b",x"73",x"b3",x"74"),
   774 => (x"4a",x"87",x"df",x"02"),
   775 => (x"fe",x"c2",x"8a",x"c2"),
   776 => (x"92",x"49",x"bf",x"e8"),
   777 => (x"bf",x"cc",x"c3",x"c3"),
   778 => (x"c3",x"80",x"72",x"48"),
   779 => (x"71",x"58",x"ec",x"c3"),
   780 => (x"c2",x"30",x"c4",x"48"),
   781 => (x"c0",x"58",x"f8",x"fe"),
   782 => (x"c3",x"c3",x"87",x"e9"),
   783 => (x"c3",x"4b",x"bf",x"d0"),
   784 => (x"c3",x"48",x"e8",x"c3"),
   785 => (x"78",x"bf",x"d4",x"c3"),
   786 => (x"bf",x"f0",x"fe",x"c2"),
   787 => (x"c2",x"87",x"c9",x"02"),
   788 => (x"49",x"bf",x"e8",x"fe"),
   789 => (x"87",x"c7",x"31",x"c4"),
   790 => (x"bf",x"d8",x"c3",x"c3"),
   791 => (x"c2",x"31",x"c4",x"49"),
   792 => (x"c3",x"59",x"f8",x"fe"),
   793 => (x"26",x"5b",x"e8",x"c3"),
   794 => (x"26",x"4b",x"26",x"4c"),
   795 => (x"5b",x"5e",x"0e",x"4f"),
   796 => (x"f0",x"0e",x"5d",x"5c"),
   797 => (x"59",x"a6",x"c8",x"86"),
   798 => (x"ff",x"ff",x"ff",x"cf"),
   799 => (x"7e",x"c0",x"4c",x"f8"),
   800 => (x"d8",x"02",x"66",x"c4"),
   801 => (x"e4",x"f6",x"c2",x"87"),
   802 => (x"c2",x"78",x"c0",x"48"),
   803 => (x"c3",x"48",x"dc",x"f6"),
   804 => (x"78",x"bf",x"e8",x"c3"),
   805 => (x"48",x"e0",x"f6",x"c2"),
   806 => (x"bf",x"e4",x"c3",x"c3"),
   807 => (x"c5",x"ff",x"c2",x"78"),
   808 => (x"c2",x"50",x"c0",x"48"),
   809 => (x"49",x"bf",x"f4",x"fe"),
   810 => (x"bf",x"e4",x"f6",x"c2"),
   811 => (x"03",x"aa",x"71",x"4a"),
   812 => (x"72",x"87",x"cc",x"c4"),
   813 => (x"05",x"99",x"cf",x"49"),
   814 => (x"c0",x"87",x"ea",x"c0"),
   815 => (x"c2",x"48",x"e8",x"f9"),
   816 => (x"78",x"bf",x"dc",x"f6"),
   817 => (x"1e",x"e8",x"f6",x"c2"),
   818 => (x"bf",x"dc",x"f6",x"c2"),
   819 => (x"dc",x"f6",x"c2",x"49"),
   820 => (x"78",x"a1",x"c1",x"48"),
   821 => (x"fd",x"df",x"ff",x"71"),
   822 => (x"c0",x"86",x"c4",x"87"),
   823 => (x"c2",x"48",x"e4",x"f9"),
   824 => (x"cc",x"78",x"e8",x"f6"),
   825 => (x"e4",x"f9",x"c0",x"87"),
   826 => (x"e0",x"c0",x"48",x"bf"),
   827 => (x"e8",x"f9",x"c0",x"80"),
   828 => (x"e4",x"f6",x"c2",x"58"),
   829 => (x"80",x"c1",x"48",x"bf"),
   830 => (x"58",x"e8",x"f6",x"c2"),
   831 => (x"00",x"0e",x"64",x"27"),
   832 => (x"bf",x"97",x"bf",x"00"),
   833 => (x"c2",x"02",x"9d",x"4d"),
   834 => (x"e5",x"c3",x"87",x"e5"),
   835 => (x"de",x"c2",x"02",x"ad"),
   836 => (x"e4",x"f9",x"c0",x"87"),
   837 => (x"a3",x"cb",x"4b",x"bf"),
   838 => (x"cf",x"4c",x"11",x"49"),
   839 => (x"d2",x"c1",x"05",x"ac"),
   840 => (x"df",x"49",x"75",x"87"),
   841 => (x"cd",x"89",x"c1",x"99"),
   842 => (x"f8",x"fe",x"c2",x"91"),
   843 => (x"4a",x"a3",x"c1",x"81"),
   844 => (x"a3",x"c3",x"51",x"12"),
   845 => (x"c5",x"51",x"12",x"4a"),
   846 => (x"51",x"12",x"4a",x"a3"),
   847 => (x"12",x"4a",x"a3",x"c7"),
   848 => (x"4a",x"a3",x"c9",x"51"),
   849 => (x"a3",x"ce",x"51",x"12"),
   850 => (x"d0",x"51",x"12",x"4a"),
   851 => (x"51",x"12",x"4a",x"a3"),
   852 => (x"12",x"4a",x"a3",x"d2"),
   853 => (x"4a",x"a3",x"d4",x"51"),
   854 => (x"a3",x"d6",x"51",x"12"),
   855 => (x"d8",x"51",x"12",x"4a"),
   856 => (x"51",x"12",x"4a",x"a3"),
   857 => (x"12",x"4a",x"a3",x"dc"),
   858 => (x"4a",x"a3",x"de",x"51"),
   859 => (x"7e",x"c1",x"51",x"12"),
   860 => (x"74",x"87",x"fc",x"c0"),
   861 => (x"05",x"99",x"c8",x"49"),
   862 => (x"74",x"87",x"ed",x"c0"),
   863 => (x"05",x"99",x"d0",x"49"),
   864 => (x"e0",x"c0",x"87",x"d3"),
   865 => (x"cc",x"c0",x"02",x"66"),
   866 => (x"c0",x"49",x"73",x"87"),
   867 => (x"70",x"0f",x"66",x"e0"),
   868 => (x"d3",x"c0",x"02",x"98"),
   869 => (x"c0",x"05",x"6e",x"87"),
   870 => (x"fe",x"c2",x"87",x"c6"),
   871 => (x"50",x"c0",x"48",x"f8"),
   872 => (x"bf",x"e4",x"f9",x"c0"),
   873 => (x"87",x"eb",x"c2",x"48"),
   874 => (x"48",x"c5",x"ff",x"c2"),
   875 => (x"c2",x"7e",x"50",x"c0"),
   876 => (x"49",x"bf",x"f4",x"fe"),
   877 => (x"bf",x"e4",x"f6",x"c2"),
   878 => (x"04",x"aa",x"71",x"4a"),
   879 => (x"cf",x"87",x"f4",x"fb"),
   880 => (x"f8",x"ff",x"ff",x"ff"),
   881 => (x"e8",x"c3",x"c3",x"4c"),
   882 => (x"c8",x"c0",x"05",x"bf"),
   883 => (x"f0",x"fe",x"c2",x"87"),
   884 => (x"fc",x"c1",x"02",x"bf"),
   885 => (x"e0",x"f6",x"c2",x"87"),
   886 => (x"c4",x"eb",x"49",x"bf"),
   887 => (x"e4",x"f6",x"c2",x"87"),
   888 => (x"48",x"a6",x"c4",x"58"),
   889 => (x"bf",x"e0",x"f6",x"c2"),
   890 => (x"f0",x"fe",x"c2",x"78"),
   891 => (x"db",x"c0",x"02",x"bf"),
   892 => (x"49",x"66",x"c4",x"87"),
   893 => (x"a9",x"74",x"99",x"74"),
   894 => (x"87",x"c8",x"c0",x"02"),
   895 => (x"c0",x"48",x"a6",x"c8"),
   896 => (x"87",x"e7",x"c0",x"78"),
   897 => (x"c1",x"48",x"a6",x"c8"),
   898 => (x"87",x"df",x"c0",x"78"),
   899 => (x"cf",x"49",x"66",x"c4"),
   900 => (x"a9",x"99",x"f8",x"ff"),
   901 => (x"87",x"c8",x"c0",x"02"),
   902 => (x"c0",x"48",x"a6",x"cc"),
   903 => (x"87",x"c5",x"c0",x"78"),
   904 => (x"c1",x"48",x"a6",x"cc"),
   905 => (x"48",x"a6",x"c8",x"78"),
   906 => (x"c8",x"78",x"66",x"cc"),
   907 => (x"e0",x"c0",x"05",x"66"),
   908 => (x"49",x"66",x"c4",x"87"),
   909 => (x"fe",x"c2",x"89",x"c2"),
   910 => (x"91",x"4a",x"bf",x"e8"),
   911 => (x"bf",x"cc",x"c3",x"c3"),
   912 => (x"dc",x"f6",x"c2",x"4a"),
   913 => (x"78",x"a1",x"72",x"48"),
   914 => (x"48",x"e4",x"f6",x"c2"),
   915 => (x"d2",x"f9",x"78",x"c0"),
   916 => (x"cf",x"48",x"c0",x"87"),
   917 => (x"f8",x"ff",x"ff",x"ff"),
   918 => (x"26",x"8e",x"f0",x"4c"),
   919 => (x"26",x"4c",x"26",x"4d"),
   920 => (x"00",x"4f",x"26",x"4b"),
   921 => (x"00",x"00",x"00",x"00"),
   922 => (x"ff",x"ff",x"ff",x"ff"),
   923 => (x"48",x"d0",x"ff",x"1e"),
   924 => (x"26",x"78",x"e0",x"c0"),
   925 => (x"e9",x"c1",x"1e",x"4f"),
   926 => (x"49",x"70",x"87",x"f7"),
   927 => (x"87",x"c6",x"02",x"99"),
   928 => (x"05",x"a9",x"fb",x"c0"),
   929 => (x"48",x"71",x"87",x"f0"),
   930 => (x"5e",x"0e",x"4f",x"26"),
   931 => (x"71",x"0e",x"5c",x"5b"),
   932 => (x"c1",x"4c",x"c0",x"4b"),
   933 => (x"70",x"87",x"da",x"e9"),
   934 => (x"c0",x"02",x"99",x"49"),
   935 => (x"ec",x"c0",x"87",x"fa"),
   936 => (x"f3",x"c0",x"02",x"a9"),
   937 => (x"a9",x"fb",x"c0",x"87"),
   938 => (x"87",x"ec",x"c0",x"02"),
   939 => (x"ac",x"b7",x"66",x"cc"),
   940 => (x"d0",x"87",x"c7",x"03"),
   941 => (x"87",x"c2",x"02",x"66"),
   942 => (x"99",x"71",x"53",x"71"),
   943 => (x"c1",x"87",x"c2",x"02"),
   944 => (x"ec",x"e8",x"c1",x"84"),
   945 => (x"99",x"49",x"70",x"87"),
   946 => (x"c0",x"87",x"cd",x"02"),
   947 => (x"c7",x"02",x"a9",x"ec"),
   948 => (x"a9",x"fb",x"c0",x"87"),
   949 => (x"87",x"d4",x"ff",x"05"),
   950 => (x"c3",x"02",x"66",x"d0"),
   951 => (x"7b",x"97",x"c0",x"87"),
   952 => (x"05",x"a9",x"fb",x"c0"),
   953 => (x"4a",x"74",x"87",x"c7"),
   954 => (x"c2",x"8a",x"0a",x"c0"),
   955 => (x"72",x"4a",x"74",x"87"),
   956 => (x"26",x"4c",x"26",x"48"),
   957 => (x"1e",x"4f",x"26",x"4b"),
   958 => (x"87",x"f5",x"e7",x"c1"),
   959 => (x"c0",x"4a",x"49",x"70"),
   960 => (x"c9",x"04",x"aa",x"f0"),
   961 => (x"aa",x"f9",x"c0",x"87"),
   962 => (x"c0",x"87",x"c3",x"01"),
   963 => (x"c1",x"c1",x"8a",x"f0"),
   964 => (x"87",x"c9",x"04",x"aa"),
   965 => (x"01",x"aa",x"da",x"c1"),
   966 => (x"f7",x"c0",x"87",x"c3"),
   967 => (x"26",x"48",x"72",x"8a"),
   968 => (x"5b",x"5e",x"0e",x"4f"),
   969 => (x"f8",x"0e",x"5d",x"5c"),
   970 => (x"c0",x"4c",x"71",x"86"),
   971 => (x"e3",x"e7",x"c1",x"7e"),
   972 => (x"c0",x"4b",x"c0",x"87"),
   973 => (x"bf",x"97",x"c4",x"ff"),
   974 => (x"04",x"a9",x"c0",x"49"),
   975 => (x"f4",x"fc",x"87",x"cf"),
   976 => (x"c0",x"83",x"c1",x"87"),
   977 => (x"bf",x"97",x"c4",x"ff"),
   978 => (x"f1",x"06",x"ab",x"49"),
   979 => (x"c4",x"ff",x"c0",x"87"),
   980 => (x"d0",x"02",x"bf",x"97"),
   981 => (x"d8",x"e6",x"c1",x"87"),
   982 => (x"99",x"49",x"70",x"87"),
   983 => (x"c0",x"87",x"c6",x"02"),
   984 => (x"f0",x"05",x"a9",x"ec"),
   985 => (x"c1",x"4b",x"c0",x"87"),
   986 => (x"70",x"87",x"c6",x"e6"),
   987 => (x"c0",x"e6",x"c1",x"4d"),
   988 => (x"58",x"a6",x"c8",x"87"),
   989 => (x"87",x"f9",x"e5",x"c1"),
   990 => (x"83",x"c1",x"4a",x"70"),
   991 => (x"97",x"49",x"a4",x"c8"),
   992 => (x"05",x"ad",x"49",x"69"),
   993 => (x"a4",x"c9",x"87",x"da"),
   994 => (x"49",x"69",x"97",x"49"),
   995 => (x"05",x"a9",x"66",x"c4"),
   996 => (x"a4",x"ca",x"87",x"ce"),
   997 => (x"49",x"69",x"97",x"49"),
   998 => (x"87",x"c4",x"05",x"aa"),
   999 => (x"87",x"d0",x"7e",x"c1"),
  1000 => (x"02",x"ad",x"ec",x"c0"),
  1001 => (x"fb",x"c0",x"87",x"c6"),
  1002 => (x"87",x"c4",x"05",x"ad"),
  1003 => (x"7e",x"c1",x"4b",x"c0"),
  1004 => (x"f2",x"fe",x"02",x"6e"),
  1005 => (x"87",x"f4",x"fa",x"87"),
  1006 => (x"8e",x"f8",x"48",x"73"),
  1007 => (x"4c",x"26",x"4d",x"26"),
  1008 => (x"4f",x"26",x"4b",x"26"),
  1009 => (x"1e",x"73",x"1e",x"00"),
  1010 => (x"c8",x"4b",x"d4",x"ff"),
  1011 => (x"d0",x"ff",x"4a",x"66"),
  1012 => (x"78",x"c5",x"c8",x"48"),
  1013 => (x"c1",x"48",x"d4",x"ff"),
  1014 => (x"7b",x"11",x"78",x"d4"),
  1015 => (x"f9",x"05",x"8a",x"c1"),
  1016 => (x"48",x"d0",x"ff",x"87"),
  1017 => (x"4b",x"26",x"78",x"c4"),
  1018 => (x"5e",x"0e",x"4f",x"26"),
  1019 => (x"0e",x"5d",x"5c",x"5b"),
  1020 => (x"7e",x"71",x"86",x"f8"),
  1021 => (x"c3",x"c3",x"1e",x"6e"),
  1022 => (x"db",x"e4",x"49",x"fc"),
  1023 => (x"70",x"86",x"c4",x"87"),
  1024 => (x"e4",x"c4",x"02",x"98"),
  1025 => (x"e4",x"e8",x"c1",x"87"),
  1026 => (x"49",x"6e",x"4c",x"bf"),
  1027 => (x"c8",x"87",x"d2",x"fc"),
  1028 => (x"98",x"70",x"58",x"a6"),
  1029 => (x"c4",x"87",x"c5",x"05"),
  1030 => (x"78",x"c1",x"48",x"a6"),
  1031 => (x"c5",x"48",x"d0",x"ff"),
  1032 => (x"48",x"d4",x"ff",x"78"),
  1033 => (x"c4",x"78",x"d5",x"c1"),
  1034 => (x"89",x"c1",x"49",x"66"),
  1035 => (x"e8",x"c1",x"31",x"c6"),
  1036 => (x"4a",x"bf",x"97",x"dc"),
  1037 => (x"ff",x"b0",x"71",x"48"),
  1038 => (x"ff",x"78",x"08",x"d4"),
  1039 => (x"78",x"c4",x"48",x"d0"),
  1040 => (x"97",x"f8",x"c3",x"c3"),
  1041 => (x"99",x"d0",x"49",x"bf"),
  1042 => (x"c5",x"87",x"dd",x"02"),
  1043 => (x"48",x"d4",x"ff",x"78"),
  1044 => (x"c0",x"78",x"d6",x"c1"),
  1045 => (x"48",x"d4",x"ff",x"4a"),
  1046 => (x"c1",x"78",x"ff",x"c3"),
  1047 => (x"aa",x"e0",x"c0",x"82"),
  1048 => (x"ff",x"87",x"f2",x"04"),
  1049 => (x"78",x"c4",x"48",x"d0"),
  1050 => (x"c3",x"48",x"d4",x"ff"),
  1051 => (x"d0",x"ff",x"78",x"ff"),
  1052 => (x"ff",x"78",x"c5",x"48"),
  1053 => (x"d3",x"c1",x"48",x"d4"),
  1054 => (x"ff",x"78",x"c1",x"78"),
  1055 => (x"78",x"c4",x"48",x"d0"),
  1056 => (x"06",x"ac",x"b7",x"c0"),
  1057 => (x"c3",x"87",x"cb",x"c2"),
  1058 => (x"4b",x"bf",x"c4",x"c4"),
  1059 => (x"73",x"7e",x"74",x"8c"),
  1060 => (x"dd",x"c1",x"02",x"9b"),
  1061 => (x"4d",x"c0",x"c8",x"87"),
  1062 => (x"ab",x"b7",x"c0",x"8b"),
  1063 => (x"c8",x"87",x"c6",x"03"),
  1064 => (x"c0",x"4d",x"a3",x"c0"),
  1065 => (x"f8",x"c3",x"c3",x"4b"),
  1066 => (x"d0",x"49",x"bf",x"97"),
  1067 => (x"87",x"cf",x"02",x"99"),
  1068 => (x"c3",x"c3",x"1e",x"c0"),
  1069 => (x"d5",x"e6",x"49",x"fc"),
  1070 => (x"70",x"86",x"c4",x"87"),
  1071 => (x"c2",x"87",x"d8",x"4c"),
  1072 => (x"c3",x"1e",x"e8",x"f6"),
  1073 => (x"e6",x"49",x"fc",x"c3"),
  1074 => (x"4c",x"70",x"87",x"c4"),
  1075 => (x"f6",x"c2",x"1e",x"75"),
  1076 => (x"f0",x"fb",x"49",x"e8"),
  1077 => (x"74",x"86",x"c8",x"87"),
  1078 => (x"87",x"c5",x"05",x"9c"),
  1079 => (x"ca",x"c1",x"48",x"c0"),
  1080 => (x"c3",x"1e",x"c1",x"87"),
  1081 => (x"e4",x"49",x"fc",x"c3"),
  1082 => (x"86",x"c4",x"87",x"d5"),
  1083 => (x"fe",x"05",x"9b",x"73"),
  1084 => (x"4c",x"6e",x"87",x"e3"),
  1085 => (x"06",x"ac",x"b7",x"c0"),
  1086 => (x"c3",x"c3",x"87",x"d1"),
  1087 => (x"78",x"c0",x"48",x"fc"),
  1088 => (x"78",x"c0",x"80",x"d0"),
  1089 => (x"c4",x"c3",x"80",x"f4"),
  1090 => (x"c0",x"78",x"bf",x"c8"),
  1091 => (x"fd",x"01",x"ac",x"b7"),
  1092 => (x"d0",x"ff",x"87",x"f5"),
  1093 => (x"ff",x"78",x"c5",x"48"),
  1094 => (x"d3",x"c1",x"48",x"d4"),
  1095 => (x"ff",x"78",x"c0",x"78"),
  1096 => (x"78",x"c4",x"48",x"d0"),
  1097 => (x"c2",x"c0",x"48",x"c1"),
  1098 => (x"f8",x"48",x"c0",x"87"),
  1099 => (x"26",x"4d",x"26",x"8e"),
  1100 => (x"26",x"4b",x"26",x"4c"),
  1101 => (x"5b",x"5e",x"0e",x"4f"),
  1102 => (x"fc",x"0e",x"5d",x"5c"),
  1103 => (x"c0",x"4d",x"71",x"86"),
  1104 => (x"04",x"ad",x"4c",x"4b"),
  1105 => (x"c0",x"87",x"e8",x"c0"),
  1106 => (x"74",x"1e",x"e1",x"fc"),
  1107 => (x"87",x"c4",x"02",x"9c"),
  1108 => (x"87",x"c2",x"4a",x"c0"),
  1109 => (x"49",x"72",x"4a",x"c1"),
  1110 => (x"c4",x"87",x"d2",x"ec"),
  1111 => (x"c1",x"7e",x"70",x"86"),
  1112 => (x"c2",x"05",x"6e",x"83"),
  1113 => (x"c1",x"4b",x"75",x"87"),
  1114 => (x"06",x"ab",x"75",x"84"),
  1115 => (x"6e",x"87",x"d8",x"ff"),
  1116 => (x"26",x"8e",x"fc",x"48"),
  1117 => (x"26",x"4c",x"26",x"4d"),
  1118 => (x"0e",x"4f",x"26",x"4b"),
  1119 => (x"5d",x"5c",x"5b",x"5e"),
  1120 => (x"71",x"86",x"fc",x"0e"),
  1121 => (x"91",x"de",x"49",x"4c"),
  1122 => (x"4d",x"dc",x"c5",x"c3"),
  1123 => (x"6d",x"97",x"85",x"71"),
  1124 => (x"87",x"dd",x"c1",x"02"),
  1125 => (x"bf",x"cc",x"c5",x"c3"),
  1126 => (x"71",x"81",x"74",x"49"),
  1127 => (x"70",x"87",x"d6",x"fe"),
  1128 => (x"02",x"98",x"48",x"7e"),
  1129 => (x"c3",x"87",x"f3",x"c0"),
  1130 => (x"70",x"4b",x"d0",x"c5"),
  1131 => (x"fe",x"49",x"cb",x"4a"),
  1132 => (x"74",x"87",x"cd",x"fd"),
  1133 => (x"c1",x"93",x"cc",x"4b"),
  1134 => (x"c4",x"83",x"e8",x"e8"),
  1135 => (x"fc",x"c7",x"c1",x"83"),
  1136 => (x"c1",x"49",x"74",x"7b"),
  1137 => (x"75",x"87",x"d5",x"c4"),
  1138 => (x"e0",x"e8",x"c1",x"7b"),
  1139 => (x"1e",x"49",x"bf",x"97"),
  1140 => (x"49",x"d0",x"c5",x"c3"),
  1141 => (x"87",x"e9",x"e5",x"c1"),
  1142 => (x"49",x"74",x"86",x"c4"),
  1143 => (x"87",x"fc",x"c3",x"c1"),
  1144 => (x"c5",x"c1",x"49",x"c0"),
  1145 => (x"c3",x"c3",x"87",x"d7"),
  1146 => (x"50",x"c0",x"48",x"f4"),
  1147 => (x"c7",x"e0",x"c0",x"49"),
  1148 => (x"26",x"8e",x"fc",x"87"),
  1149 => (x"26",x"4c",x"26",x"4d"),
  1150 => (x"00",x"4f",x"26",x"4b"),
  1151 => (x"64",x"61",x"6f",x"4c"),
  1152 => (x"2e",x"67",x"6e",x"69"),
  1153 => (x"00",x"00",x"2e",x"2e"),
  1154 => (x"61",x"42",x"20",x"80"),
  1155 => (x"00",x"00",x"6b",x"63"),
  1156 => (x"64",x"61",x"6f",x"4c"),
  1157 => (x"20",x"2e",x"2a",x"20"),
  1158 => (x"00",x"00",x"00",x"00"),
  1159 => (x"00",x"00",x"20",x"3a"),
  1160 => (x"61",x"42",x"20",x"80"),
  1161 => (x"00",x"00",x"6b",x"63"),
  1162 => (x"78",x"45",x"20",x"80"),
  1163 => (x"00",x"00",x"74",x"69"),
  1164 => (x"49",x"20",x"44",x"53"),
  1165 => (x"2e",x"74",x"69",x"6e"),
  1166 => (x"00",x"00",x"00",x"2e"),
  1167 => (x"00",x"00",x"4b",x"4f"),
  1168 => (x"54",x"4f",x"4f",x"42"),
  1169 => (x"20",x"20",x"20",x"20"),
  1170 => (x"00",x"4d",x"4f",x"52"),
  1171 => (x"71",x"1e",x"73",x"1e"),
  1172 => (x"c5",x"c3",x"49",x"4b"),
  1173 => (x"71",x"81",x"bf",x"cc"),
  1174 => (x"70",x"87",x"da",x"fb"),
  1175 => (x"c4",x"02",x"9a",x"4a"),
  1176 => (x"c2",x"e6",x"49",x"87"),
  1177 => (x"cc",x"c5",x"c3",x"87"),
  1178 => (x"73",x"78",x"c0",x"48"),
  1179 => (x"87",x"fa",x"c1",x"49"),
  1180 => (x"4f",x"26",x"4b",x"26"),
  1181 => (x"71",x"1e",x"73",x"1e"),
  1182 => (x"4a",x"a3",x"c4",x"4b"),
  1183 => (x"87",x"d0",x"c1",x"02"),
  1184 => (x"dc",x"02",x"8a",x"c1"),
  1185 => (x"c0",x"02",x"8a",x"87"),
  1186 => (x"05",x"8a",x"87",x"f2"),
  1187 => (x"c3",x"87",x"d3",x"c1"),
  1188 => (x"02",x"bf",x"cc",x"c5"),
  1189 => (x"48",x"87",x"cb",x"c1"),
  1190 => (x"c5",x"c3",x"88",x"c1"),
  1191 => (x"c1",x"c1",x"58",x"d0"),
  1192 => (x"cc",x"c5",x"c3",x"87"),
  1193 => (x"89",x"c6",x"49",x"bf"),
  1194 => (x"59",x"d0",x"c5",x"c3"),
  1195 => (x"03",x"a9",x"b7",x"c0"),
  1196 => (x"c3",x"87",x"ef",x"c0"),
  1197 => (x"c0",x"48",x"cc",x"c5"),
  1198 => (x"87",x"e6",x"c0",x"78"),
  1199 => (x"bf",x"c8",x"c5",x"c3"),
  1200 => (x"c3",x"87",x"df",x"02"),
  1201 => (x"48",x"bf",x"cc",x"c5"),
  1202 => (x"c5",x"c3",x"80",x"c1"),
  1203 => (x"87",x"d2",x"58",x"d0"),
  1204 => (x"bf",x"c8",x"c5",x"c3"),
  1205 => (x"c3",x"87",x"cb",x"02"),
  1206 => (x"48",x"bf",x"cc",x"c5"),
  1207 => (x"c5",x"c3",x"80",x"c6"),
  1208 => (x"49",x"73",x"58",x"d0"),
  1209 => (x"4b",x"26",x"87",x"c4"),
  1210 => (x"5e",x"0e",x"4f",x"26"),
  1211 => (x"0e",x"5d",x"5c",x"5b"),
  1212 => (x"a6",x"d0",x"86",x"f0"),
  1213 => (x"e8",x"f6",x"c2",x"59"),
  1214 => (x"c3",x"4c",x"c0",x"4d"),
  1215 => (x"c1",x"48",x"c8",x"c5"),
  1216 => (x"48",x"a6",x"c4",x"78"),
  1217 => (x"7e",x"75",x"78",x"c0"),
  1218 => (x"bf",x"cc",x"c5",x"c3"),
  1219 => (x"06",x"a8",x"c0",x"48"),
  1220 => (x"75",x"87",x"fa",x"c0"),
  1221 => (x"e8",x"f6",x"c2",x"7e"),
  1222 => (x"c0",x"02",x"98",x"48"),
  1223 => (x"fc",x"c0",x"87",x"ef"),
  1224 => (x"66",x"c8",x"1e",x"e1"),
  1225 => (x"c0",x"87",x"c4",x"02"),
  1226 => (x"c1",x"87",x"c2",x"4d"),
  1227 => (x"e4",x"49",x"75",x"4d"),
  1228 => (x"86",x"c4",x"87",x"fb"),
  1229 => (x"84",x"c1",x"7e",x"70"),
  1230 => (x"c1",x"48",x"66",x"c4"),
  1231 => (x"58",x"a6",x"c8",x"80"),
  1232 => (x"bf",x"cc",x"c5",x"c3"),
  1233 => (x"87",x"c5",x"03",x"ac"),
  1234 => (x"d1",x"ff",x"05",x"6e"),
  1235 => (x"c0",x"4d",x"6e",x"87"),
  1236 => (x"02",x"9d",x"75",x"4c"),
  1237 => (x"c0",x"87",x"e0",x"c3"),
  1238 => (x"c8",x"1e",x"e1",x"fc"),
  1239 => (x"87",x"c7",x"02",x"66"),
  1240 => (x"c0",x"48",x"a6",x"cc"),
  1241 => (x"cc",x"87",x"c5",x"78"),
  1242 => (x"78",x"c1",x"48",x"a6"),
  1243 => (x"e3",x"49",x"66",x"cc"),
  1244 => (x"86",x"c4",x"87",x"fb"),
  1245 => (x"98",x"48",x"7e",x"70"),
  1246 => (x"87",x"e8",x"c2",x"02"),
  1247 => (x"97",x"81",x"cb",x"49"),
  1248 => (x"99",x"d0",x"49",x"69"),
  1249 => (x"87",x"d6",x"c1",x"02"),
  1250 => (x"4a",x"cc",x"c9",x"c1"),
  1251 => (x"91",x"cc",x"49",x"74"),
  1252 => (x"81",x"e8",x"e8",x"c1"),
  1253 => (x"81",x"c8",x"79",x"72"),
  1254 => (x"74",x"51",x"ff",x"c3"),
  1255 => (x"c3",x"91",x"de",x"49"),
  1256 => (x"71",x"4d",x"dc",x"c5"),
  1257 => (x"97",x"c1",x"c2",x"85"),
  1258 => (x"49",x"a5",x"c1",x"7d"),
  1259 => (x"c2",x"51",x"e0",x"c0"),
  1260 => (x"bf",x"97",x"f8",x"fe"),
  1261 => (x"c1",x"87",x"d2",x"02"),
  1262 => (x"4b",x"a5",x"c2",x"84"),
  1263 => (x"4a",x"f8",x"fe",x"c2"),
  1264 => (x"f4",x"fe",x"49",x"db"),
  1265 => (x"db",x"c1",x"87",x"fa"),
  1266 => (x"49",x"a5",x"cd",x"87"),
  1267 => (x"84",x"c1",x"51",x"c0"),
  1268 => (x"6e",x"4b",x"a5",x"c2"),
  1269 => (x"fe",x"49",x"cb",x"4a"),
  1270 => (x"c1",x"87",x"e5",x"f4"),
  1271 => (x"c5",x"c1",x"87",x"c6"),
  1272 => (x"49",x"74",x"4a",x"fb"),
  1273 => (x"e8",x"c1",x"91",x"cc"),
  1274 => (x"79",x"72",x"81",x"e8"),
  1275 => (x"97",x"f8",x"fe",x"c2"),
  1276 => (x"87",x"d8",x"02",x"bf"),
  1277 => (x"91",x"de",x"49",x"74"),
  1278 => (x"c5",x"c3",x"84",x"c1"),
  1279 => (x"83",x"71",x"4b",x"dc"),
  1280 => (x"4a",x"f8",x"fe",x"c2"),
  1281 => (x"f3",x"fe",x"49",x"dd"),
  1282 => (x"87",x"d8",x"87",x"f6"),
  1283 => (x"93",x"de",x"4b",x"74"),
  1284 => (x"83",x"dc",x"c5",x"c3"),
  1285 => (x"c0",x"49",x"a3",x"cb"),
  1286 => (x"73",x"84",x"c1",x"51"),
  1287 => (x"49",x"cb",x"4a",x"6e"),
  1288 => (x"87",x"dc",x"f3",x"fe"),
  1289 => (x"c1",x"48",x"66",x"c4"),
  1290 => (x"58",x"a6",x"c8",x"80"),
  1291 => (x"c0",x"03",x"ac",x"c7"),
  1292 => (x"05",x"6e",x"87",x"c5"),
  1293 => (x"c7",x"87",x"e0",x"fc"),
  1294 => (x"e6",x"c0",x"03",x"ac"),
  1295 => (x"c8",x"c5",x"c3",x"87"),
  1296 => (x"c1",x"78",x"c0",x"48"),
  1297 => (x"74",x"4a",x"fb",x"c5"),
  1298 => (x"c1",x"91",x"cc",x"49"),
  1299 => (x"72",x"81",x"e8",x"e8"),
  1300 => (x"de",x"49",x"74",x"79"),
  1301 => (x"dc",x"c5",x"c3",x"91"),
  1302 => (x"c1",x"51",x"c0",x"81"),
  1303 => (x"04",x"ac",x"c7",x"84"),
  1304 => (x"c1",x"87",x"da",x"ff"),
  1305 => (x"c0",x"48",x"c4",x"ea"),
  1306 => (x"c1",x"80",x"f7",x"50"),
  1307 => (x"c1",x"40",x"d1",x"d3"),
  1308 => (x"c8",x"78",x"c8",x"c8"),
  1309 => (x"f4",x"c9",x"c1",x"80"),
  1310 => (x"49",x"66",x"cc",x"78"),
  1311 => (x"87",x"dc",x"f9",x"c0"),
  1312 => (x"4d",x"26",x"8e",x"f0"),
  1313 => (x"4b",x"26",x"4c",x"26"),
  1314 => (x"73",x"1e",x"4f",x"26"),
  1315 => (x"49",x"4b",x"71",x"1e"),
  1316 => (x"e8",x"c1",x"91",x"cc"),
  1317 => (x"a1",x"c8",x"81",x"e8"),
  1318 => (x"dc",x"e8",x"c1",x"4a"),
  1319 => (x"c9",x"50",x"12",x"48"),
  1320 => (x"ff",x"c0",x"4a",x"a1"),
  1321 => (x"50",x"12",x"48",x"c4"),
  1322 => (x"e8",x"c1",x"81",x"ca"),
  1323 => (x"50",x"11",x"48",x"e0"),
  1324 => (x"97",x"e0",x"e8",x"c1"),
  1325 => (x"c0",x"1e",x"49",x"bf"),
  1326 => (x"c4",x"da",x"c1",x"49"),
  1327 => (x"f8",x"49",x"73",x"87"),
  1328 => (x"8e",x"fc",x"87",x"e8"),
  1329 => (x"4f",x"26",x"4b",x"26"),
  1330 => (x"c0",x"49",x"c0",x"1e"),
  1331 => (x"26",x"87",x"ee",x"f9"),
  1332 => (x"4a",x"71",x"1e",x"4f"),
  1333 => (x"c1",x"91",x"cc",x"49"),
  1334 => (x"c8",x"81",x"e8",x"e8"),
  1335 => (x"f4",x"c3",x"c3",x"81"),
  1336 => (x"c0",x"50",x"11",x"48"),
  1337 => (x"fe",x"49",x"a2",x"f0"),
  1338 => (x"c0",x"87",x"e1",x"ee"),
  1339 => (x"87",x"c8",x"d4",x"49"),
  1340 => (x"5e",x"0e",x"4f",x"26"),
  1341 => (x"0e",x"5d",x"5c",x"5b"),
  1342 => (x"4d",x"71",x"86",x"f4"),
  1343 => (x"c1",x"91",x"cc",x"49"),
  1344 => (x"c8",x"81",x"e8",x"e8"),
  1345 => (x"a1",x"ca",x"4a",x"a1"),
  1346 => (x"48",x"a6",x"c4",x"7e"),
  1347 => (x"bf",x"f0",x"c3",x"c3"),
  1348 => (x"bf",x"97",x"6e",x"78"),
  1349 => (x"4c",x"66",x"c4",x"4b"),
  1350 => (x"48",x"12",x"2c",x"73"),
  1351 => (x"70",x"58",x"a6",x"cc"),
  1352 => (x"c9",x"84",x"c1",x"9c"),
  1353 => (x"49",x"69",x"97",x"81"),
  1354 => (x"c2",x"04",x"ac",x"b7"),
  1355 => (x"6e",x"4c",x"c0",x"87"),
  1356 => (x"c8",x"4a",x"bf",x"97"),
  1357 => (x"31",x"72",x"49",x"66"),
  1358 => (x"66",x"c4",x"b9",x"ff"),
  1359 => (x"72",x"48",x"74",x"99"),
  1360 => (x"b1",x"4a",x"70",x"30"),
  1361 => (x"59",x"f4",x"c3",x"c3"),
  1362 => (x"f8",x"cd",x"c1",x"71"),
  1363 => (x"c3",x"1e",x"c7",x"87"),
  1364 => (x"1e",x"bf",x"c4",x"c5"),
  1365 => (x"1e",x"e8",x"e8",x"c1"),
  1366 => (x"97",x"f4",x"c3",x"c3"),
  1367 => (x"e2",x"c1",x"49",x"bf"),
  1368 => (x"c0",x"49",x"75",x"87"),
  1369 => (x"e8",x"87",x"f5",x"f5"),
  1370 => (x"26",x"4d",x"26",x"8e"),
  1371 => (x"26",x"4b",x"26",x"4c"),
  1372 => (x"1e",x"73",x"1e",x"4f"),
  1373 => (x"a3",x"c2",x"4b",x"71"),
  1374 => (x"87",x"d6",x"02",x"4a"),
  1375 => (x"c0",x"05",x"8a",x"c1"),
  1376 => (x"c5",x"c3",x"87",x"e2"),
  1377 => (x"db",x"02",x"bf",x"c4"),
  1378 => (x"88",x"c1",x"48",x"87"),
  1379 => (x"58",x"c8",x"c5",x"c3"),
  1380 => (x"c5",x"c3",x"87",x"d2"),
  1381 => (x"cb",x"02",x"bf",x"c8"),
  1382 => (x"c4",x"c5",x"c3",x"87"),
  1383 => (x"80",x"c1",x"48",x"bf"),
  1384 => (x"58",x"c8",x"c5",x"c3"),
  1385 => (x"c5",x"c3",x"1e",x"c7"),
  1386 => (x"c1",x"1e",x"bf",x"c4"),
  1387 => (x"c3",x"1e",x"e8",x"e8"),
  1388 => (x"bf",x"97",x"f4",x"c3"),
  1389 => (x"73",x"87",x"cc",x"49"),
  1390 => (x"df",x"f4",x"c0",x"49"),
  1391 => (x"26",x"8e",x"f4",x"87"),
  1392 => (x"0e",x"4f",x"26",x"4b"),
  1393 => (x"5d",x"5c",x"5b",x"5e"),
  1394 => (x"86",x"cc",x"ff",x"0e"),
  1395 => (x"59",x"a6",x"e8",x"c0"),
  1396 => (x"c0",x"48",x"a6",x"cc"),
  1397 => (x"c0",x"80",x"c4",x"78"),
  1398 => (x"c0",x"80",x"c4",x"78"),
  1399 => (x"c1",x"80",x"c4",x"78"),
  1400 => (x"c4",x"78",x"66",x"c8"),
  1401 => (x"c4",x"78",x"c1",x"80"),
  1402 => (x"c3",x"78",x"c1",x"80"),
  1403 => (x"c1",x"48",x"c8",x"c5"),
  1404 => (x"df",x"cc",x"c1",x"78"),
  1405 => (x"87",x"fd",x"e1",x"87"),
  1406 => (x"87",x"f5",x"cb",x"c1"),
  1407 => (x"fb",x"c0",x"4d",x"70"),
  1408 => (x"f2",x"c1",x"02",x"ad"),
  1409 => (x"66",x"e4",x"c0",x"87"),
  1410 => (x"87",x"e7",x"c1",x"05"),
  1411 => (x"4a",x"66",x"c4",x"c1"),
  1412 => (x"7e",x"6a",x"82",x"c4"),
  1413 => (x"48",x"d0",x"c8",x"c1"),
  1414 => (x"41",x"20",x"49",x"6e"),
  1415 => (x"51",x"10",x"41",x"20"),
  1416 => (x"48",x"66",x"c4",x"c1"),
  1417 => (x"78",x"ca",x"d2",x"c1"),
  1418 => (x"81",x"c7",x"49",x"6a"),
  1419 => (x"c4",x"c1",x"51",x"75"),
  1420 => (x"81",x"c8",x"49",x"66"),
  1421 => (x"a6",x"dc",x"51",x"c1"),
  1422 => (x"c1",x"78",x"c2",x"48"),
  1423 => (x"c9",x"49",x"66",x"c4"),
  1424 => (x"c1",x"51",x"c0",x"81"),
  1425 => (x"ca",x"49",x"66",x"c4"),
  1426 => (x"c1",x"51",x"c0",x"81"),
  1427 => (x"6a",x"1e",x"d8",x"1e"),
  1428 => (x"e0",x"81",x"c8",x"49"),
  1429 => (x"86",x"c8",x"87",x"f4"),
  1430 => (x"48",x"66",x"c8",x"c1"),
  1431 => (x"c7",x"01",x"a8",x"c0"),
  1432 => (x"48",x"a6",x"d4",x"87"),
  1433 => (x"87",x"cf",x"78",x"c1"),
  1434 => (x"48",x"66",x"c8",x"c1"),
  1435 => (x"a6",x"dc",x"88",x"c1"),
  1436 => (x"ff",x"87",x"c4",x"58"),
  1437 => (x"75",x"87",x"fe",x"df"),
  1438 => (x"f3",x"cb",x"02",x"9d"),
  1439 => (x"48",x"66",x"d4",x"87"),
  1440 => (x"a8",x"66",x"cc",x"c1"),
  1441 => (x"87",x"e8",x"cb",x"03"),
  1442 => (x"c9",x"c1",x"7e",x"c0"),
  1443 => (x"4d",x"70",x"87",x"e3"),
  1444 => (x"88",x"c6",x"c1",x"48"),
  1445 => (x"70",x"58",x"a6",x"c8"),
  1446 => (x"d6",x"c1",x"02",x"98"),
  1447 => (x"88",x"c9",x"48",x"87"),
  1448 => (x"70",x"58",x"a6",x"c8"),
  1449 => (x"d9",x"c5",x"02",x"98"),
  1450 => (x"88",x"c1",x"48",x"87"),
  1451 => (x"70",x"58",x"a6",x"c8"),
  1452 => (x"f8",x"c2",x"02",x"98"),
  1453 => (x"88",x"c3",x"48",x"87"),
  1454 => (x"70",x"58",x"a6",x"c8"),
  1455 => (x"87",x"cf",x"02",x"98"),
  1456 => (x"c8",x"88",x"c1",x"48"),
  1457 => (x"98",x"70",x"58",x"a6"),
  1458 => (x"87",x"f6",x"c4",x"02"),
  1459 => (x"c0",x"87",x"c0",x"ca"),
  1460 => (x"c8",x"c1",x"7e",x"f0"),
  1461 => (x"4d",x"70",x"87",x"db"),
  1462 => (x"02",x"ad",x"ec",x"c0"),
  1463 => (x"7e",x"75",x"87",x"c2"),
  1464 => (x"02",x"ad",x"ec",x"c0"),
  1465 => (x"c8",x"c1",x"87",x"cd"),
  1466 => (x"4d",x"70",x"87",x"c7"),
  1467 => (x"05",x"ad",x"ec",x"c0"),
  1468 => (x"c0",x"87",x"f3",x"ff"),
  1469 => (x"c1",x"05",x"66",x"e4"),
  1470 => (x"ec",x"c0",x"87",x"ea"),
  1471 => (x"87",x"c4",x"02",x"ad"),
  1472 => (x"87",x"ed",x"c7",x"c1"),
  1473 => (x"1e",x"ca",x"1e",x"c0"),
  1474 => (x"cc",x"4b",x"66",x"dc"),
  1475 => (x"66",x"cc",x"c1",x"93"),
  1476 => (x"4c",x"a3",x"c4",x"83"),
  1477 => (x"dd",x"ff",x"49",x"6c"),
  1478 => (x"1e",x"c1",x"87",x"f0"),
  1479 => (x"49",x"6c",x"1e",x"de"),
  1480 => (x"87",x"e6",x"dd",x"ff"),
  1481 => (x"d2",x"c1",x"86",x"d0"),
  1482 => (x"a3",x"c8",x"7b",x"ca"),
  1483 => (x"51",x"66",x"dc",x"49"),
  1484 => (x"c0",x"49",x"a3",x"c9"),
  1485 => (x"ca",x"51",x"66",x"e0"),
  1486 => (x"51",x"6e",x"49",x"a3"),
  1487 => (x"c1",x"48",x"66",x"dc"),
  1488 => (x"a6",x"e0",x"c0",x"80"),
  1489 => (x"48",x"66",x"d4",x"58"),
  1490 => (x"04",x"a8",x"66",x"d8"),
  1491 => (x"66",x"d4",x"87",x"cb"),
  1492 => (x"d8",x"80",x"c1",x"48"),
  1493 => (x"fc",x"c7",x"58",x"a6"),
  1494 => (x"48",x"66",x"d8",x"87"),
  1495 => (x"a6",x"dc",x"88",x"c1"),
  1496 => (x"87",x"f1",x"c7",x"58"),
  1497 => (x"87",x"cd",x"dc",x"ff"),
  1498 => (x"e8",x"c7",x"4d",x"70"),
  1499 => (x"c6",x"de",x"ff",x"87"),
  1500 => (x"58",x"a6",x"d0",x"87"),
  1501 => (x"06",x"a8",x"66",x"d0"),
  1502 => (x"d0",x"87",x"c6",x"c0"),
  1503 => (x"66",x"cc",x"48",x"a6"),
  1504 => (x"f2",x"dd",x"ff",x"78"),
  1505 => (x"a8",x"ec",x"c0",x"87"),
  1506 => (x"87",x"f6",x"c1",x"05"),
  1507 => (x"05",x"66",x"e4",x"c0"),
  1508 => (x"d4",x"87",x"e6",x"c1"),
  1509 => (x"91",x"cc",x"49",x"66"),
  1510 => (x"81",x"66",x"c4",x"c1"),
  1511 => (x"6a",x"4a",x"a1",x"c4"),
  1512 => (x"4a",x"a1",x"c8",x"4c"),
  1513 => (x"c1",x"52",x"66",x"cc"),
  1514 => (x"c1",x"79",x"d1",x"d3"),
  1515 => (x"70",x"87",x"c2",x"c5"),
  1516 => (x"db",x"02",x"9d",x"4d"),
  1517 => (x"ad",x"fb",x"c0",x"87"),
  1518 => (x"87",x"d4",x"c0",x"02"),
  1519 => (x"c4",x"c1",x"54",x"75"),
  1520 => (x"4d",x"70",x"87",x"ef"),
  1521 => (x"c7",x"c0",x"02",x"9d"),
  1522 => (x"ad",x"fb",x"c0",x"87"),
  1523 => (x"87",x"ec",x"ff",x"05"),
  1524 => (x"c2",x"54",x"e0",x"c0"),
  1525 => (x"97",x"c0",x"54",x"c1"),
  1526 => (x"48",x"66",x"d4",x"7c"),
  1527 => (x"04",x"a8",x"66",x"d8"),
  1528 => (x"d4",x"87",x"cb",x"c0"),
  1529 => (x"80",x"c1",x"48",x"66"),
  1530 => (x"c5",x"58",x"a6",x"d8"),
  1531 => (x"66",x"d8",x"87",x"e7"),
  1532 => (x"dc",x"88",x"c1",x"48"),
  1533 => (x"dc",x"c5",x"58",x"a6"),
  1534 => (x"f8",x"d9",x"ff",x"87"),
  1535 => (x"c5",x"4d",x"70",x"87"),
  1536 => (x"66",x"cc",x"87",x"d3"),
  1537 => (x"66",x"e4",x"c0",x"48"),
  1538 => (x"f4",x"c4",x"05",x"a8"),
  1539 => (x"a6",x"e8",x"c0",x"87"),
  1540 => (x"ff",x"78",x"c0",x"48"),
  1541 => (x"70",x"87",x"e0",x"db"),
  1542 => (x"da",x"db",x"ff",x"7e"),
  1543 => (x"a6",x"f0",x"c0",x"87"),
  1544 => (x"a8",x"ec",x"c0",x"58"),
  1545 => (x"87",x"c7",x"c0",x"05"),
  1546 => (x"78",x"6e",x"48",x"a6"),
  1547 => (x"c1",x"87",x"c4",x"c0"),
  1548 => (x"d4",x"87",x"fe",x"c2"),
  1549 => (x"91",x"cc",x"49",x"66"),
  1550 => (x"48",x"66",x"c4",x"c1"),
  1551 => (x"a6",x"c8",x"80",x"71"),
  1552 => (x"4a",x"66",x"c4",x"58"),
  1553 => (x"66",x"c4",x"82",x"c8"),
  1554 => (x"6e",x"81",x"ca",x"49"),
  1555 => (x"66",x"ec",x"c0",x"51"),
  1556 => (x"6e",x"81",x"c1",x"49"),
  1557 => (x"71",x"48",x"c1",x"89"),
  1558 => (x"c1",x"49",x"70",x"30"),
  1559 => (x"7a",x"97",x"71",x"89"),
  1560 => (x"bf",x"f0",x"c3",x"c3"),
  1561 => (x"97",x"29",x"6e",x"49"),
  1562 => (x"71",x"48",x"4a",x"6a"),
  1563 => (x"a6",x"f4",x"c0",x"98"),
  1564 => (x"48",x"66",x"c4",x"58"),
  1565 => (x"a6",x"cc",x"80",x"c4"),
  1566 => (x"bf",x"66",x"c8",x"58"),
  1567 => (x"66",x"e4",x"c0",x"4c"),
  1568 => (x"a8",x"66",x"cc",x"48"),
  1569 => (x"87",x"c5",x"c0",x"02"),
  1570 => (x"c2",x"c0",x"7e",x"c0"),
  1571 => (x"6e",x"7e",x"c1",x"87"),
  1572 => (x"1e",x"e0",x"c0",x"1e"),
  1573 => (x"d7",x"ff",x"49",x"74"),
  1574 => (x"86",x"c8",x"87",x"f0"),
  1575 => (x"b7",x"c0",x"4d",x"70"),
  1576 => (x"d4",x"c1",x"06",x"ad"),
  1577 => (x"c8",x"84",x"75",x"87"),
  1578 => (x"c0",x"49",x"bf",x"66"),
  1579 => (x"89",x"74",x"81",x"e0"),
  1580 => (x"dc",x"c8",x"c1",x"4b"),
  1581 => (x"e1",x"fe",x"71",x"4a"),
  1582 => (x"84",x"c2",x"87",x"c6"),
  1583 => (x"e8",x"c0",x"7e",x"74"),
  1584 => (x"80",x"c1",x"48",x"66"),
  1585 => (x"58",x"a6",x"ec",x"c0"),
  1586 => (x"49",x"66",x"f0",x"c0"),
  1587 => (x"a9",x"70",x"81",x"c1"),
  1588 => (x"87",x"c5",x"c0",x"02"),
  1589 => (x"c2",x"c0",x"4c",x"c0"),
  1590 => (x"74",x"4c",x"c1",x"87"),
  1591 => (x"bf",x"66",x"cc",x"1e"),
  1592 => (x"81",x"e0",x"c0",x"49"),
  1593 => (x"71",x"89",x"66",x"c4"),
  1594 => (x"49",x"66",x"c8",x"1e"),
  1595 => (x"87",x"da",x"d6",x"ff"),
  1596 => (x"b7",x"c0",x"86",x"c8"),
  1597 => (x"c5",x"ff",x"01",x"a8"),
  1598 => (x"66",x"e8",x"c0",x"87"),
  1599 => (x"87",x"d3",x"c0",x"02"),
  1600 => (x"c9",x"49",x"66",x"c4"),
  1601 => (x"66",x"e8",x"c0",x"81"),
  1602 => (x"48",x"66",x"c4",x"51"),
  1603 => (x"78",x"f2",x"d3",x"c1"),
  1604 => (x"c4",x"87",x"ce",x"c0"),
  1605 => (x"81",x"c9",x"49",x"66"),
  1606 => (x"66",x"c4",x"51",x"c2"),
  1607 => (x"e3",x"eb",x"c2",x"48"),
  1608 => (x"48",x"66",x"d4",x"78"),
  1609 => (x"04",x"a8",x"66",x"d8"),
  1610 => (x"d4",x"87",x"cb",x"c0"),
  1611 => (x"80",x"c1",x"48",x"66"),
  1612 => (x"c0",x"58",x"a6",x"d8"),
  1613 => (x"66",x"d8",x"87",x"d1"),
  1614 => (x"dc",x"88",x"c1",x"48"),
  1615 => (x"c6",x"c0",x"58",x"a6"),
  1616 => (x"f0",x"d4",x"ff",x"87"),
  1617 => (x"cc",x"4d",x"70",x"87"),
  1618 => (x"78",x"c0",x"48",x"a6"),
  1619 => (x"ff",x"87",x"c6",x"c0"),
  1620 => (x"70",x"87",x"e2",x"d4"),
  1621 => (x"66",x"e0",x"c0",x"4d"),
  1622 => (x"c0",x"80",x"c1",x"48"),
  1623 => (x"75",x"58",x"a6",x"e4"),
  1624 => (x"cb",x"c0",x"02",x"9d"),
  1625 => (x"48",x"66",x"d4",x"87"),
  1626 => (x"a8",x"66",x"cc",x"c1"),
  1627 => (x"87",x"d8",x"f4",x"04"),
  1628 => (x"c7",x"48",x"66",x"d4"),
  1629 => (x"e1",x"c0",x"03",x"a8"),
  1630 => (x"4c",x"66",x"d4",x"87"),
  1631 => (x"48",x"c8",x"c5",x"c3"),
  1632 => (x"49",x"74",x"78",x"c0"),
  1633 => (x"c4",x"c1",x"91",x"cc"),
  1634 => (x"a1",x"c4",x"81",x"66"),
  1635 => (x"c0",x"4a",x"6a",x"4a"),
  1636 => (x"84",x"c1",x"79",x"52"),
  1637 => (x"ff",x"04",x"ac",x"c7"),
  1638 => (x"e4",x"c0",x"87",x"e2"),
  1639 => (x"e2",x"c0",x"02",x"66"),
  1640 => (x"66",x"c4",x"c1",x"87"),
  1641 => (x"81",x"d4",x"c1",x"49"),
  1642 => (x"4a",x"66",x"c4",x"c1"),
  1643 => (x"c0",x"82",x"dc",x"c1"),
  1644 => (x"d1",x"d3",x"c1",x"52"),
  1645 => (x"66",x"c4",x"c1",x"79"),
  1646 => (x"81",x"d8",x"c1",x"49"),
  1647 => (x"79",x"e0",x"c8",x"c1"),
  1648 => (x"c1",x"87",x"d6",x"c0"),
  1649 => (x"c1",x"49",x"66",x"c4"),
  1650 => (x"c4",x"c1",x"81",x"d4"),
  1651 => (x"d8",x"c1",x"4a",x"66"),
  1652 => (x"e8",x"c8",x"c1",x"82"),
  1653 => (x"c8",x"d3",x"c1",x"7a"),
  1654 => (x"f1",x"d5",x"c1",x"79"),
  1655 => (x"66",x"c4",x"c1",x"4a"),
  1656 => (x"81",x"e0",x"c1",x"49"),
  1657 => (x"d2",x"ff",x"79",x"72"),
  1658 => (x"66",x"d0",x"87",x"c2"),
  1659 => (x"8e",x"cc",x"ff",x"48"),
  1660 => (x"4c",x"26",x"4d",x"26"),
  1661 => (x"4f",x"26",x"4b",x"26"),
  1662 => (x"c3",x"1e",x"c7",x"1e"),
  1663 => (x"1e",x"bf",x"c4",x"c5"),
  1664 => (x"1e",x"e8",x"e8",x"c1"),
  1665 => (x"97",x"f4",x"c3",x"c3"),
  1666 => (x"f6",x"ee",x"49",x"bf"),
  1667 => (x"e8",x"e8",x"c1",x"87"),
  1668 => (x"d5",x"e4",x"c0",x"49"),
  1669 => (x"26",x"8e",x"f4",x"87"),
  1670 => (x"00",x"00",x"00",x"4f"),
  1671 => (x"00",x"00",x"00",x"00"),
  1672 => (x"00",x"00",x"00",x"00"),
  1673 => (x"00",x"00",x"00",x"01"),
  1674 => (x"00",x"00",x"11",x"7b"),
  1675 => (x"00",x"00",x"31",x"5c"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"00",x"00",x"11",x"7b"),
  1678 => (x"00",x"00",x"31",x"7a"),
  1679 => (x"00",x"00",x"00",x"00"),
  1680 => (x"00",x"00",x"11",x"7b"),
  1681 => (x"00",x"00",x"31",x"98"),
  1682 => (x"00",x"00",x"00",x"00"),
  1683 => (x"00",x"00",x"11",x"7b"),
  1684 => (x"00",x"00",x"31",x"b6"),
  1685 => (x"00",x"00",x"00",x"00"),
  1686 => (x"00",x"00",x"11",x"7b"),
  1687 => (x"00",x"00",x"31",x"d4"),
  1688 => (x"00",x"00",x"00",x"00"),
  1689 => (x"00",x"00",x"11",x"7b"),
  1690 => (x"00",x"00",x"31",x"f2"),
  1691 => (x"00",x"00",x"00",x"00"),
  1692 => (x"00",x"00",x"11",x"7b"),
  1693 => (x"00",x"00",x"32",x"10"),
  1694 => (x"00",x"00",x"00",x"00"),
  1695 => (x"00",x"00",x"14",x"d1"),
  1696 => (x"00",x"00",x"00",x"00"),
  1697 => (x"00",x"00",x"00",x"00"),
  1698 => (x"00",x"00",x"12",x"74"),
  1699 => (x"00",x"00",x"00",x"00"),
  1700 => (x"00",x"00",x"00",x"00"),
  1701 => (x"00",x"00",x"12",x"40"),
  1702 => (x"db",x"86",x"fc",x"1e"),
  1703 => (x"fc",x"7e",x"70",x"87"),
  1704 => (x"1e",x"4f",x"26",x"8e"),
  1705 => (x"c0",x"48",x"f0",x"fe"),
  1706 => (x"79",x"09",x"cd",x"78"),
  1707 => (x"1e",x"4f",x"26",x"09"),
  1708 => (x"49",x"d8",x"ea",x"c1"),
  1709 => (x"4f",x"26",x"87",x"ed"),
  1710 => (x"bf",x"f0",x"fe",x"1e"),
  1711 => (x"1e",x"4f",x"26",x"48"),
  1712 => (x"c1",x"48",x"f0",x"fe"),
  1713 => (x"1e",x"4f",x"26",x"78"),
  1714 => (x"c0",x"48",x"f0",x"fe"),
  1715 => (x"1e",x"4f",x"26",x"78"),
  1716 => (x"97",x"c0",x"4a",x"71"),
  1717 => (x"49",x"a2",x"c1",x"7a"),
  1718 => (x"a2",x"ca",x"51",x"c0"),
  1719 => (x"cb",x"51",x"c0",x"49"),
  1720 => (x"51",x"c0",x"49",x"a2"),
  1721 => (x"5e",x"0e",x"4f",x"26"),
  1722 => (x"f0",x"0e",x"5c",x"5b"),
  1723 => (x"ca",x"4c",x"71",x"86"),
  1724 => (x"69",x"97",x"49",x"a4"),
  1725 => (x"4b",x"a4",x"cb",x"7e"),
  1726 => (x"c8",x"48",x"6b",x"97"),
  1727 => (x"80",x"c1",x"58",x"a6"),
  1728 => (x"c7",x"58",x"a6",x"cc"),
  1729 => (x"58",x"a6",x"d0",x"98"),
  1730 => (x"66",x"cc",x"48",x"6e"),
  1731 => (x"87",x"db",x"05",x"a8"),
  1732 => (x"97",x"7e",x"69",x"97"),
  1733 => (x"a6",x"c8",x"48",x"6b"),
  1734 => (x"cc",x"80",x"c1",x"58"),
  1735 => (x"98",x"c7",x"58",x"a6"),
  1736 => (x"6e",x"58",x"a6",x"d0"),
  1737 => (x"a8",x"66",x"cc",x"48"),
  1738 => (x"fe",x"87",x"e5",x"02"),
  1739 => (x"a4",x"cc",x"87",x"d9"),
  1740 => (x"49",x"6b",x"97",x"4a"),
  1741 => (x"dc",x"49",x"a1",x"72"),
  1742 => (x"6b",x"97",x"51",x"66"),
  1743 => (x"c1",x"48",x"6e",x"7e"),
  1744 => (x"58",x"a6",x"c8",x"80"),
  1745 => (x"a6",x"cc",x"98",x"c7"),
  1746 => (x"7b",x"97",x"70",x"58"),
  1747 => (x"fd",x"87",x"de",x"c1"),
  1748 => (x"8e",x"f0",x"87",x"ed"),
  1749 => (x"4b",x"26",x"4c",x"26"),
  1750 => (x"5e",x"0e",x"4f",x"26"),
  1751 => (x"0e",x"5d",x"5c",x"5b"),
  1752 => (x"4d",x"71",x"86",x"f4"),
  1753 => (x"c1",x"7e",x"6d",x"97"),
  1754 => (x"6c",x"97",x"4c",x"a5"),
  1755 => (x"58",x"a6",x"c8",x"48"),
  1756 => (x"66",x"c4",x"48",x"6e"),
  1757 => (x"87",x"c5",x"05",x"a8"),
  1758 => (x"e6",x"c0",x"48",x"ff"),
  1759 => (x"87",x"c7",x"fd",x"87"),
  1760 => (x"97",x"49",x"a5",x"c2"),
  1761 => (x"a3",x"71",x"4b",x"6c"),
  1762 => (x"4b",x"6b",x"97",x"4b"),
  1763 => (x"6e",x"7e",x"6c",x"97"),
  1764 => (x"c8",x"80",x"c1",x"48"),
  1765 => (x"98",x"c7",x"58",x"a6"),
  1766 => (x"70",x"58",x"a6",x"cc"),
  1767 => (x"de",x"fc",x"7c",x"97"),
  1768 => (x"f4",x"48",x"73",x"87"),
  1769 => (x"26",x"4d",x"26",x"8e"),
  1770 => (x"26",x"4b",x"26",x"4c"),
  1771 => (x"5b",x"5e",x"0e",x"4f"),
  1772 => (x"86",x"f4",x"0e",x"5c"),
  1773 => (x"e0",x"87",x"d0",x"fc"),
  1774 => (x"c0",x"49",x"4c",x"bf"),
  1775 => (x"02",x"99",x"c0",x"e0"),
  1776 => (x"74",x"87",x"ea",x"c0"),
  1777 => (x"9a",x"ff",x"c3",x"4a"),
  1778 => (x"97",x"c4",x"c9",x"c3"),
  1779 => (x"c9",x"c3",x"49",x"bf"),
  1780 => (x"51",x"72",x"81",x"c6"),
  1781 => (x"97",x"c4",x"c9",x"c3"),
  1782 => (x"48",x"6e",x"7e",x"bf"),
  1783 => (x"a6",x"c8",x"80",x"c1"),
  1784 => (x"cc",x"98",x"c7",x"58"),
  1785 => (x"c9",x"c3",x"58",x"a6"),
  1786 => (x"66",x"c8",x"48",x"c4"),
  1787 => (x"d0",x"49",x"74",x"50"),
  1788 => (x"c1",x"02",x"99",x"c0"),
  1789 => (x"c9",x"c3",x"87",x"c0"),
  1790 => (x"7e",x"bf",x"97",x"ce"),
  1791 => (x"97",x"cf",x"c9",x"c3"),
  1792 => (x"a6",x"c8",x"48",x"bf"),
  1793 => (x"c4",x"48",x"6e",x"58"),
  1794 => (x"c0",x"02",x"a8",x"66"),
  1795 => (x"c9",x"c3",x"87",x"e8"),
  1796 => (x"49",x"bf",x"97",x"ce"),
  1797 => (x"81",x"d0",x"c9",x"c3"),
  1798 => (x"08",x"e0",x"48",x"11"),
  1799 => (x"ce",x"c9",x"c3",x"78"),
  1800 => (x"6e",x"7e",x"bf",x"97"),
  1801 => (x"c8",x"80",x"c1",x"48"),
  1802 => (x"98",x"c7",x"58",x"a6"),
  1803 => (x"c3",x"58",x"a6",x"cc"),
  1804 => (x"c8",x"48",x"ce",x"c9"),
  1805 => (x"bf",x"e4",x"50",x"66"),
  1806 => (x"e0",x"c0",x"49",x"4b"),
  1807 => (x"c0",x"02",x"99",x"c0"),
  1808 => (x"4a",x"73",x"87",x"ea"),
  1809 => (x"c3",x"9a",x"ff",x"c3"),
  1810 => (x"bf",x"97",x"d8",x"c9"),
  1811 => (x"da",x"c9",x"c3",x"49"),
  1812 => (x"c3",x"51",x"72",x"81"),
  1813 => (x"bf",x"97",x"d8",x"c9"),
  1814 => (x"c1",x"48",x"6e",x"7e"),
  1815 => (x"58",x"a6",x"c8",x"80"),
  1816 => (x"a6",x"cc",x"98",x"c7"),
  1817 => (x"d8",x"c9",x"c3",x"58"),
  1818 => (x"50",x"66",x"c8",x"48"),
  1819 => (x"c0",x"d0",x"49",x"73"),
  1820 => (x"c0",x"c1",x"02",x"99"),
  1821 => (x"e2",x"c9",x"c3",x"87"),
  1822 => (x"c3",x"7e",x"bf",x"97"),
  1823 => (x"bf",x"97",x"e3",x"c9"),
  1824 => (x"58",x"a6",x"c8",x"48"),
  1825 => (x"66",x"c4",x"48",x"6e"),
  1826 => (x"e8",x"c0",x"02",x"a8"),
  1827 => (x"e2",x"c9",x"c3",x"87"),
  1828 => (x"c3",x"49",x"bf",x"97"),
  1829 => (x"11",x"81",x"e4",x"c9"),
  1830 => (x"78",x"08",x"e4",x"48"),
  1831 => (x"97",x"e2",x"c9",x"c3"),
  1832 => (x"48",x"6e",x"7e",x"bf"),
  1833 => (x"a6",x"c8",x"80",x"c1"),
  1834 => (x"cc",x"98",x"c7",x"58"),
  1835 => (x"c9",x"c3",x"58",x"a6"),
  1836 => (x"66",x"c8",x"48",x"e2"),
  1837 => (x"87",x"c0",x"f8",x"50"),
  1838 => (x"c2",x"f8",x"7e",x"70"),
  1839 => (x"26",x"8e",x"f4",x"87"),
  1840 => (x"26",x"4b",x"26",x"4c"),
  1841 => (x"c9",x"c3",x"1e",x"4f"),
  1842 => (x"c2",x"f8",x"49",x"c4"),
  1843 => (x"d8",x"c9",x"c3",x"87"),
  1844 => (x"87",x"fb",x"f7",x"49"),
  1845 => (x"49",x"ed",x"ee",x"c1"),
  1846 => (x"c3",x"87",x"c8",x"f7"),
  1847 => (x"4f",x"26",x"87",x"f2"),
  1848 => (x"c3",x"1e",x"73",x"1e"),
  1849 => (x"f9",x"49",x"c4",x"c9"),
  1850 => (x"4a",x"70",x"87",x"f0"),
  1851 => (x"04",x"aa",x"b7",x"c0"),
  1852 => (x"c3",x"87",x"cc",x"c2"),
  1853 => (x"c9",x"05",x"aa",x"f0"),
  1854 => (x"c8",x"f6",x"c1",x"87"),
  1855 => (x"c1",x"78",x"c1",x"48"),
  1856 => (x"e0",x"c3",x"87",x"ed"),
  1857 => (x"87",x"c9",x"05",x"aa"),
  1858 => (x"48",x"cc",x"f6",x"c1"),
  1859 => (x"de",x"c1",x"78",x"c1"),
  1860 => (x"cc",x"f6",x"c1",x"87"),
  1861 => (x"87",x"c6",x"02",x"bf"),
  1862 => (x"4b",x"a2",x"c0",x"c2"),
  1863 => (x"4b",x"72",x"87",x"c2"),
  1864 => (x"bf",x"c8",x"f6",x"c1"),
  1865 => (x"87",x"e0",x"c0",x"02"),
  1866 => (x"b7",x"c4",x"49",x"73"),
  1867 => (x"f6",x"c1",x"91",x"29"),
  1868 => (x"4a",x"73",x"81",x"d0"),
  1869 => (x"92",x"c2",x"9a",x"cf"),
  1870 => (x"30",x"72",x"48",x"c1"),
  1871 => (x"ba",x"ff",x"4a",x"70"),
  1872 => (x"98",x"69",x"48",x"72"),
  1873 => (x"87",x"db",x"79",x"70"),
  1874 => (x"b7",x"c4",x"49",x"73"),
  1875 => (x"f6",x"c1",x"91",x"29"),
  1876 => (x"4a",x"73",x"81",x"d0"),
  1877 => (x"92",x"c2",x"9a",x"cf"),
  1878 => (x"30",x"72",x"48",x"c3"),
  1879 => (x"69",x"48",x"4a",x"70"),
  1880 => (x"c1",x"79",x"70",x"b0"),
  1881 => (x"c0",x"48",x"cc",x"f6"),
  1882 => (x"c8",x"f6",x"c1",x"78"),
  1883 => (x"c3",x"78",x"c0",x"48"),
  1884 => (x"f7",x"49",x"c4",x"c9"),
  1885 => (x"4a",x"70",x"87",x"e4"),
  1886 => (x"03",x"aa",x"b7",x"c0"),
  1887 => (x"c0",x"87",x"f4",x"fd"),
  1888 => (x"26",x"4b",x"26",x"48"),
  1889 => (x"00",x"00",x"00",x"4f"),
  1890 => (x"00",x"00",x"00",x"00"),
  1891 => (x"00",x"00",x"00",x"00"),
  1892 => (x"00",x"00",x"00",x"00"),
  1893 => (x"00",x"00",x"00",x"00"),
  1894 => (x"00",x"00",x"00",x"00"),
  1895 => (x"00",x"00",x"00",x"00"),
  1896 => (x"00",x"00",x"00",x"00"),
  1897 => (x"00",x"00",x"00",x"00"),
  1898 => (x"00",x"00",x"00",x"00"),
  1899 => (x"00",x"00",x"00",x"00"),
  1900 => (x"00",x"00",x"00",x"00"),
  1901 => (x"00",x"00",x"00",x"00"),
  1902 => (x"00",x"00",x"00",x"00"),
  1903 => (x"00",x"00",x"00",x"00"),
  1904 => (x"00",x"00",x"00",x"00"),
  1905 => (x"00",x"00",x"00",x"00"),
  1906 => (x"00",x"00",x"00",x"00"),
  1907 => (x"00",x"00",x"00",x"00"),
  1908 => (x"72",x"4a",x"c0",x"1e"),
  1909 => (x"c1",x"91",x"c4",x"49"),
  1910 => (x"c0",x"81",x"d0",x"f6"),
  1911 => (x"d0",x"82",x"c1",x"79"),
  1912 => (x"ee",x"04",x"aa",x"b7"),
  1913 => (x"0e",x"4f",x"26",x"87"),
  1914 => (x"5d",x"5c",x"5b",x"5e"),
  1915 => (x"f3",x"4d",x"71",x"0e"),
  1916 => (x"4a",x"75",x"87",x"d5"),
  1917 => (x"92",x"2a",x"b7",x"c4"),
  1918 => (x"82",x"d0",x"f6",x"c1"),
  1919 => (x"9c",x"cf",x"4c",x"75"),
  1920 => (x"49",x"6a",x"94",x"c2"),
  1921 => (x"c3",x"2b",x"74",x"4b"),
  1922 => (x"74",x"48",x"c2",x"9b"),
  1923 => (x"ff",x"4c",x"70",x"30"),
  1924 => (x"71",x"48",x"74",x"bc"),
  1925 => (x"f2",x"7a",x"70",x"98"),
  1926 => (x"48",x"73",x"87",x"e5"),
  1927 => (x"4c",x"26",x"4d",x"26"),
  1928 => (x"4f",x"26",x"4b",x"26"),
  1929 => (x"48",x"d0",x"ff",x"1e"),
  1930 => (x"71",x"78",x"e1",x"c8"),
  1931 => (x"08",x"d4",x"ff",x"48"),
  1932 => (x"1e",x"4f",x"26",x"78"),
  1933 => (x"c8",x"48",x"d0",x"ff"),
  1934 => (x"48",x"71",x"78",x"e1"),
  1935 => (x"78",x"08",x"d4",x"ff"),
  1936 => (x"ff",x"48",x"66",x"c4"),
  1937 => (x"26",x"78",x"08",x"d4"),
  1938 => (x"4a",x"71",x"1e",x"4f"),
  1939 => (x"1e",x"49",x"66",x"c4"),
  1940 => (x"de",x"ff",x"49",x"72"),
  1941 => (x"48",x"d0",x"ff",x"87"),
  1942 => (x"fc",x"78",x"e0",x"c0"),
  1943 => (x"1e",x"4f",x"26",x"8e"),
  1944 => (x"4a",x"71",x"1e",x"73"),
  1945 => (x"ab",x"b7",x"c2",x"4b"),
  1946 => (x"a3",x"87",x"c8",x"03"),
  1947 => (x"ff",x"c3",x"4a",x"49"),
  1948 => (x"ce",x"87",x"c7",x"9a"),
  1949 => (x"c3",x"4a",x"49",x"a3"),
  1950 => (x"66",x"c8",x"9a",x"ff"),
  1951 => (x"49",x"72",x"1e",x"49"),
  1952 => (x"fc",x"87",x"c6",x"ff"),
  1953 => (x"26",x"4b",x"26",x"8e"),
  1954 => (x"d0",x"ff",x"1e",x"4f"),
  1955 => (x"78",x"c9",x"c8",x"48"),
  1956 => (x"d4",x"ff",x"48",x"71"),
  1957 => (x"4f",x"26",x"78",x"08"),
  1958 => (x"49",x"4a",x"71",x"1e"),
  1959 => (x"d0",x"ff",x"87",x"eb"),
  1960 => (x"26",x"78",x"c8",x"48"),
  1961 => (x"1e",x"73",x"1e",x"4f"),
  1962 => (x"c9",x"c3",x"4b",x"71"),
  1963 => (x"c3",x"02",x"bf",x"f8"),
  1964 => (x"87",x"eb",x"c2",x"87"),
  1965 => (x"c8",x"48",x"d0",x"ff"),
  1966 => (x"48",x"73",x"78",x"c9"),
  1967 => (x"ff",x"b0",x"e0",x"c0"),
  1968 => (x"c3",x"78",x"08",x"d4"),
  1969 => (x"c0",x"48",x"ec",x"c9"),
  1970 => (x"02",x"66",x"c8",x"78"),
  1971 => (x"ff",x"c3",x"87",x"c5"),
  1972 => (x"c0",x"87",x"c2",x"49"),
  1973 => (x"f4",x"c9",x"c3",x"49"),
  1974 => (x"02",x"66",x"cc",x"59"),
  1975 => (x"d5",x"c5",x"87",x"c6"),
  1976 => (x"87",x"c4",x"4a",x"d5"),
  1977 => (x"4a",x"ff",x"ff",x"cf"),
  1978 => (x"5a",x"f8",x"c9",x"c3"),
  1979 => (x"48",x"f8",x"c9",x"c3"),
  1980 => (x"4b",x"26",x"78",x"c1"),
  1981 => (x"5e",x"0e",x"4f",x"26"),
  1982 => (x"0e",x"5d",x"5c",x"5b"),
  1983 => (x"c9",x"c3",x"4d",x"71"),
  1984 => (x"75",x"4b",x"bf",x"f4"),
  1985 => (x"87",x"cb",x"02",x"9d"),
  1986 => (x"c1",x"91",x"c8",x"49"),
  1987 => (x"71",x"4a",x"dc",x"fa"),
  1988 => (x"c1",x"87",x"c4",x"82"),
  1989 => (x"c0",x"4a",x"dc",x"fe"),
  1990 => (x"73",x"49",x"12",x"4c"),
  1991 => (x"f0",x"c9",x"c3",x"99"),
  1992 => (x"b8",x"71",x"48",x"bf"),
  1993 => (x"78",x"08",x"d4",x"ff"),
  1994 => (x"84",x"2b",x"b7",x"c1"),
  1995 => (x"04",x"ac",x"b7",x"c8"),
  1996 => (x"c9",x"c3",x"87",x"e7"),
  1997 => (x"c8",x"48",x"bf",x"ec"),
  1998 => (x"f0",x"c9",x"c3",x"80"),
  1999 => (x"26",x"4d",x"26",x"58"),
  2000 => (x"26",x"4b",x"26",x"4c"),
  2001 => (x"1e",x"73",x"1e",x"4f"),
  2002 => (x"4a",x"13",x"4b",x"71"),
  2003 => (x"87",x"cb",x"02",x"9a"),
  2004 => (x"e1",x"fe",x"49",x"72"),
  2005 => (x"9a",x"4a",x"13",x"87"),
  2006 => (x"26",x"87",x"f5",x"05"),
  2007 => (x"1e",x"4f",x"26",x"4b"),
  2008 => (x"bf",x"ec",x"c9",x"c3"),
  2009 => (x"ec",x"c9",x"c3",x"49"),
  2010 => (x"78",x"a1",x"c1",x"48"),
  2011 => (x"a9",x"b7",x"c0",x"c4"),
  2012 => (x"ff",x"87",x"db",x"03"),
  2013 => (x"c9",x"c3",x"48",x"d4"),
  2014 => (x"c3",x"78",x"bf",x"f0"),
  2015 => (x"49",x"bf",x"ec",x"c9"),
  2016 => (x"48",x"ec",x"c9",x"c3"),
  2017 => (x"c4",x"78",x"a1",x"c1"),
  2018 => (x"04",x"a9",x"b7",x"c0"),
  2019 => (x"d0",x"ff",x"87",x"e5"),
  2020 => (x"c3",x"78",x"c8",x"48"),
  2021 => (x"c0",x"48",x"f8",x"c9"),
  2022 => (x"00",x"4f",x"26",x"78"),
  2023 => (x"00",x"00",x"00",x"00"),
  2024 => (x"00",x"00",x"00",x"00"),
  2025 => (x"5f",x"00",x"00",x"00"),
  2026 => (x"00",x"00",x"00",x"5f"),
  2027 => (x"00",x"03",x"03",x"00"),
  2028 => (x"00",x"00",x"03",x"03"),
  2029 => (x"14",x"7f",x"7f",x"14"),
  2030 => (x"00",x"14",x"7f",x"7f"),
  2031 => (x"6b",x"2e",x"24",x"00"),
  2032 => (x"00",x"12",x"3a",x"6b"),
  2033 => (x"18",x"36",x"6a",x"4c"),
  2034 => (x"00",x"32",x"56",x"6c"),
  2035 => (x"59",x"4f",x"7e",x"30"),
  2036 => (x"40",x"68",x"3a",x"77"),
  2037 => (x"07",x"04",x"00",x"00"),
  2038 => (x"00",x"00",x"00",x"03"),
  2039 => (x"3e",x"1c",x"00",x"00"),
  2040 => (x"00",x"00",x"41",x"63"),
  2041 => (x"63",x"41",x"00",x"00"),
  2042 => (x"00",x"00",x"1c",x"3e"),
  2043 => (x"1c",x"3e",x"2a",x"08"),
  2044 => (x"08",x"2a",x"3e",x"1c"),
  2045 => (x"3e",x"08",x"08",x"00"),
  2046 => (x"00",x"08",x"08",x"3e"),
  2047 => (x"e0",x"80",x"00",x"00"),
  2048 => (x"00",x"00",x"00",x"60"),
  2049 => (x"08",x"08",x"08",x"00"),
  2050 => (x"00",x"08",x"08",x"08"),
  2051 => (x"60",x"00",x"00",x"00"),
  2052 => (x"00",x"00",x"00",x"60"),
  2053 => (x"18",x"30",x"60",x"40"),
  2054 => (x"01",x"03",x"06",x"0c"),
  2055 => (x"59",x"7f",x"3e",x"00"),
  2056 => (x"00",x"3e",x"7f",x"4d"),
  2057 => (x"7f",x"06",x"04",x"00"),
  2058 => (x"00",x"00",x"00",x"7f"),
  2059 => (x"71",x"63",x"42",x"00"),
  2060 => (x"00",x"46",x"4f",x"59"),
  2061 => (x"49",x"63",x"22",x"00"),
  2062 => (x"00",x"36",x"7f",x"49"),
  2063 => (x"13",x"16",x"1c",x"18"),
  2064 => (x"00",x"10",x"7f",x"7f"),
  2065 => (x"45",x"67",x"27",x"00"),
  2066 => (x"00",x"39",x"7d",x"45"),
  2067 => (x"4b",x"7e",x"3c",x"00"),
  2068 => (x"00",x"30",x"79",x"49"),
  2069 => (x"71",x"01",x"01",x"00"),
  2070 => (x"00",x"07",x"0f",x"79"),
  2071 => (x"49",x"7f",x"36",x"00"),
  2072 => (x"00",x"36",x"7f",x"49"),
  2073 => (x"49",x"4f",x"06",x"00"),
  2074 => (x"00",x"1e",x"3f",x"69"),
  2075 => (x"66",x"00",x"00",x"00"),
  2076 => (x"00",x"00",x"00",x"66"),
  2077 => (x"e6",x"80",x"00",x"00"),
  2078 => (x"00",x"00",x"00",x"66"),
  2079 => (x"14",x"08",x"08",x"00"),
  2080 => (x"00",x"22",x"22",x"14"),
  2081 => (x"14",x"14",x"14",x"00"),
  2082 => (x"00",x"14",x"14",x"14"),
  2083 => (x"14",x"22",x"22",x"00"),
  2084 => (x"00",x"08",x"08",x"14"),
  2085 => (x"51",x"03",x"02",x"00"),
  2086 => (x"00",x"06",x"0f",x"59"),
  2087 => (x"5d",x"41",x"7f",x"3e"),
  2088 => (x"00",x"1e",x"1f",x"55"),
  2089 => (x"09",x"7f",x"7e",x"00"),
  2090 => (x"00",x"7e",x"7f",x"09"),
  2091 => (x"49",x"7f",x"7f",x"00"),
  2092 => (x"00",x"36",x"7f",x"49"),
  2093 => (x"63",x"3e",x"1c",x"00"),
  2094 => (x"00",x"41",x"41",x"41"),
  2095 => (x"41",x"7f",x"7f",x"00"),
  2096 => (x"00",x"1c",x"3e",x"63"),
  2097 => (x"49",x"7f",x"7f",x"00"),
  2098 => (x"00",x"41",x"41",x"49"),
  2099 => (x"09",x"7f",x"7f",x"00"),
  2100 => (x"00",x"01",x"01",x"09"),
  2101 => (x"41",x"7f",x"3e",x"00"),
  2102 => (x"00",x"7a",x"7b",x"49"),
  2103 => (x"08",x"7f",x"7f",x"00"),
  2104 => (x"00",x"7f",x"7f",x"08"),
  2105 => (x"7f",x"41",x"00",x"00"),
  2106 => (x"00",x"00",x"41",x"7f"),
  2107 => (x"40",x"60",x"20",x"00"),
  2108 => (x"00",x"3f",x"7f",x"40"),
  2109 => (x"1c",x"08",x"7f",x"7f"),
  2110 => (x"00",x"41",x"63",x"36"),
  2111 => (x"40",x"7f",x"7f",x"00"),
  2112 => (x"00",x"40",x"40",x"40"),
  2113 => (x"0c",x"06",x"7f",x"7f"),
  2114 => (x"00",x"7f",x"7f",x"06"),
  2115 => (x"0c",x"06",x"7f",x"7f"),
  2116 => (x"00",x"7f",x"7f",x"18"),
  2117 => (x"41",x"7f",x"3e",x"00"),
  2118 => (x"00",x"3e",x"7f",x"41"),
  2119 => (x"09",x"7f",x"7f",x"00"),
  2120 => (x"00",x"06",x"0f",x"09"),
  2121 => (x"61",x"41",x"7f",x"3e"),
  2122 => (x"00",x"40",x"7e",x"7f"),
  2123 => (x"09",x"7f",x"7f",x"00"),
  2124 => (x"00",x"66",x"7f",x"19"),
  2125 => (x"4d",x"6f",x"26",x"00"),
  2126 => (x"00",x"32",x"7b",x"59"),
  2127 => (x"7f",x"01",x"01",x"00"),
  2128 => (x"00",x"01",x"01",x"7f"),
  2129 => (x"40",x"7f",x"3f",x"00"),
  2130 => (x"00",x"3f",x"7f",x"40"),
  2131 => (x"70",x"3f",x"0f",x"00"),
  2132 => (x"00",x"0f",x"3f",x"70"),
  2133 => (x"18",x"30",x"7f",x"7f"),
  2134 => (x"00",x"7f",x"7f",x"30"),
  2135 => (x"1c",x"36",x"63",x"41"),
  2136 => (x"41",x"63",x"36",x"1c"),
  2137 => (x"7c",x"06",x"03",x"01"),
  2138 => (x"01",x"03",x"06",x"7c"),
  2139 => (x"4d",x"59",x"71",x"61"),
  2140 => (x"00",x"41",x"43",x"47"),
  2141 => (x"7f",x"7f",x"00",x"00"),
  2142 => (x"00",x"00",x"41",x"41"),
  2143 => (x"0c",x"06",x"03",x"01"),
  2144 => (x"40",x"60",x"30",x"18"),
  2145 => (x"41",x"41",x"00",x"00"),
  2146 => (x"00",x"00",x"7f",x"7f"),
  2147 => (x"03",x"06",x"0c",x"08"),
  2148 => (x"00",x"08",x"0c",x"06"),
  2149 => (x"80",x"80",x"80",x"80"),
  2150 => (x"00",x"80",x"80",x"80"),
  2151 => (x"03",x"00",x"00",x"00"),
  2152 => (x"00",x"00",x"04",x"07"),
  2153 => (x"54",x"74",x"20",x"00"),
  2154 => (x"00",x"78",x"7c",x"54"),
  2155 => (x"44",x"7f",x"7f",x"00"),
  2156 => (x"00",x"38",x"7c",x"44"),
  2157 => (x"44",x"7c",x"38",x"00"),
  2158 => (x"00",x"00",x"44",x"44"),
  2159 => (x"44",x"7c",x"38",x"00"),
  2160 => (x"00",x"7f",x"7f",x"44"),
  2161 => (x"54",x"7c",x"38",x"00"),
  2162 => (x"00",x"18",x"5c",x"54"),
  2163 => (x"7f",x"7e",x"04",x"00"),
  2164 => (x"00",x"00",x"05",x"05"),
  2165 => (x"a4",x"bc",x"18",x"00"),
  2166 => (x"00",x"7c",x"fc",x"a4"),
  2167 => (x"04",x"7f",x"7f",x"00"),
  2168 => (x"00",x"78",x"7c",x"04"),
  2169 => (x"3d",x"00",x"00",x"00"),
  2170 => (x"00",x"00",x"40",x"7d"),
  2171 => (x"80",x"80",x"80",x"00"),
  2172 => (x"00",x"00",x"7d",x"fd"),
  2173 => (x"10",x"7f",x"7f",x"00"),
  2174 => (x"00",x"44",x"6c",x"38"),
  2175 => (x"3f",x"00",x"00",x"00"),
  2176 => (x"00",x"00",x"40",x"7f"),
  2177 => (x"18",x"0c",x"7c",x"7c"),
  2178 => (x"00",x"78",x"7c",x"0c"),
  2179 => (x"04",x"7c",x"7c",x"00"),
  2180 => (x"00",x"78",x"7c",x"04"),
  2181 => (x"44",x"7c",x"38",x"00"),
  2182 => (x"00",x"38",x"7c",x"44"),
  2183 => (x"24",x"fc",x"fc",x"00"),
  2184 => (x"00",x"18",x"3c",x"24"),
  2185 => (x"24",x"3c",x"18",x"00"),
  2186 => (x"00",x"fc",x"fc",x"24"),
  2187 => (x"04",x"7c",x"7c",x"00"),
  2188 => (x"00",x"08",x"0c",x"04"),
  2189 => (x"54",x"5c",x"48",x"00"),
  2190 => (x"00",x"20",x"74",x"54"),
  2191 => (x"7f",x"3f",x"04",x"00"),
  2192 => (x"00",x"00",x"44",x"44"),
  2193 => (x"40",x"7c",x"3c",x"00"),
  2194 => (x"00",x"7c",x"7c",x"40"),
  2195 => (x"60",x"3c",x"1c",x"00"),
  2196 => (x"00",x"1c",x"3c",x"60"),
  2197 => (x"30",x"60",x"7c",x"3c"),
  2198 => (x"00",x"3c",x"7c",x"60"),
  2199 => (x"10",x"38",x"6c",x"44"),
  2200 => (x"00",x"44",x"6c",x"38"),
  2201 => (x"e0",x"bc",x"1c",x"00"),
  2202 => (x"00",x"1c",x"3c",x"60"),
  2203 => (x"74",x"64",x"44",x"00"),
  2204 => (x"00",x"44",x"4c",x"5c"),
  2205 => (x"3e",x"08",x"08",x"00"),
  2206 => (x"00",x"41",x"41",x"77"),
  2207 => (x"7f",x"00",x"00",x"00"),
  2208 => (x"00",x"00",x"00",x"7f"),
  2209 => (x"77",x"41",x"41",x"00"),
  2210 => (x"00",x"08",x"08",x"3e"),
  2211 => (x"03",x"01",x"01",x"02"),
  2212 => (x"00",x"01",x"02",x"02"),
  2213 => (x"7f",x"7f",x"7f",x"7f"),
  2214 => (x"00",x"7f",x"7f",x"7f"),
  2215 => (x"1c",x"1c",x"08",x"08"),
  2216 => (x"7f",x"7f",x"3e",x"3e"),
  2217 => (x"3e",x"3e",x"7f",x"7f"),
  2218 => (x"08",x"08",x"1c",x"1c"),
  2219 => (x"7c",x"18",x"10",x"00"),
  2220 => (x"00",x"10",x"18",x"7c"),
  2221 => (x"7c",x"30",x"10",x"00"),
  2222 => (x"00",x"10",x"30",x"7c"),
  2223 => (x"60",x"60",x"30",x"10"),
  2224 => (x"00",x"06",x"1e",x"78"),
  2225 => (x"18",x"3c",x"66",x"42"),
  2226 => (x"00",x"42",x"66",x"3c"),
  2227 => (x"c2",x"6a",x"38",x"78"),
  2228 => (x"00",x"38",x"6c",x"c6"),
  2229 => (x"60",x"00",x"00",x"60"),
  2230 => (x"00",x"60",x"00",x"00"),
  2231 => (x"5c",x"5b",x"5e",x"0e"),
  2232 => (x"86",x"fc",x"0e",x"5d"),
  2233 => (x"ca",x"c3",x"7e",x"71"),
  2234 => (x"c0",x"4c",x"bf",x"c0"),
  2235 => (x"c4",x"1e",x"c0",x"4b"),
  2236 => (x"c4",x"02",x"ab",x"66"),
  2237 => (x"c2",x"4d",x"c0",x"87"),
  2238 => (x"75",x"4d",x"c1",x"87"),
  2239 => (x"ee",x"49",x"73",x"1e"),
  2240 => (x"86",x"c8",x"87",x"e3"),
  2241 => (x"ef",x"49",x"e0",x"c0"),
  2242 => (x"a4",x"c4",x"87",x"ec"),
  2243 => (x"f0",x"49",x"6a",x"4a"),
  2244 => (x"ca",x"f1",x"87",x"f3"),
  2245 => (x"c1",x"84",x"cc",x"87"),
  2246 => (x"ab",x"b7",x"c8",x"83"),
  2247 => (x"87",x"cd",x"ff",x"04"),
  2248 => (x"4d",x"26",x"8e",x"fc"),
  2249 => (x"4b",x"26",x"4c",x"26"),
  2250 => (x"71",x"1e",x"4f",x"26"),
  2251 => (x"c4",x"ca",x"c3",x"4a"),
  2252 => (x"c4",x"ca",x"c3",x"5a"),
  2253 => (x"49",x"78",x"c7",x"48"),
  2254 => (x"26",x"87",x"e1",x"fe"),
  2255 => (x"1e",x"73",x"1e",x"4f"),
  2256 => (x"0b",x"fc",x"4b",x"71"),
  2257 => (x"4a",x"73",x"0b",x"7b"),
  2258 => (x"c0",x"c1",x"9a",x"c1"),
  2259 => (x"c7",x"ed",x"49",x"a2"),
  2260 => (x"d0",x"da",x"c2",x"87"),
  2261 => (x"26",x"4b",x"26",x"5b"),
  2262 => (x"4a",x"71",x"1e",x"4f"),
  2263 => (x"72",x"1e",x"66",x"c4"),
  2264 => (x"87",x"fb",x"eb",x"49"),
  2265 => (x"4f",x"26",x"8e",x"fc"),
  2266 => (x"48",x"d4",x"ff",x"1e"),
  2267 => (x"ff",x"78",x"ff",x"c3"),
  2268 => (x"e1",x"c0",x"48",x"d0"),
  2269 => (x"48",x"d4",x"ff",x"78"),
  2270 => (x"48",x"71",x"78",x"c1"),
  2271 => (x"d4",x"ff",x"30",x"c4"),
  2272 => (x"d0",x"ff",x"78",x"08"),
  2273 => (x"78",x"e0",x"c0",x"48"),
  2274 => (x"5e",x"0e",x"4f",x"26"),
  2275 => (x"0e",x"5d",x"5c",x"5b"),
  2276 => (x"7e",x"c0",x"86",x"f4"),
  2277 => (x"ec",x"48",x"a6",x"c8"),
  2278 => (x"80",x"fc",x"78",x"bf"),
  2279 => (x"bf",x"c0",x"ca",x"c3"),
  2280 => (x"c8",x"ca",x"c3",x"78"),
  2281 => (x"bf",x"e8",x"4c",x"bf"),
  2282 => (x"cc",x"da",x"c2",x"4d"),
  2283 => (x"ef",x"e4",x"49",x"bf"),
  2284 => (x"e8",x"49",x"c7",x"87"),
  2285 => (x"49",x"70",x"87",x"f1"),
  2286 => (x"d0",x"05",x"99",x"c2"),
  2287 => (x"c4",x"da",x"c2",x"87"),
  2288 => (x"b9",x"ff",x"49",x"bf"),
  2289 => (x"c1",x"99",x"66",x"c8"),
  2290 => (x"f9",x"c1",x"02",x"99"),
  2291 => (x"49",x"e8",x"cf",x"87"),
  2292 => (x"70",x"87",x"fd",x"ca"),
  2293 => (x"e8",x"49",x"c7",x"4b"),
  2294 => (x"98",x"70",x"87",x"cd"),
  2295 => (x"c8",x"87",x"c9",x"05"),
  2296 => (x"99",x"c1",x"49",x"66"),
  2297 => (x"87",x"fe",x"c0",x"02"),
  2298 => (x"ec",x"48",x"a6",x"c8"),
  2299 => (x"ef",x"e3",x"78",x"bf"),
  2300 => (x"ca",x"49",x"73",x"87"),
  2301 => (x"98",x"70",x"87",x"e6"),
  2302 => (x"c2",x"87",x"d7",x"02"),
  2303 => (x"49",x"bf",x"c0",x"da"),
  2304 => (x"da",x"c2",x"b9",x"c1"),
  2305 => (x"fd",x"71",x"59",x"c4"),
  2306 => (x"e8",x"cf",x"87",x"de"),
  2307 => (x"87",x"c0",x"ca",x"49"),
  2308 => (x"49",x"c7",x"4b",x"70"),
  2309 => (x"70",x"87",x"d0",x"e7"),
  2310 => (x"cb",x"ff",x"05",x"98"),
  2311 => (x"49",x"66",x"c8",x"87"),
  2312 => (x"ff",x"05",x"99",x"c1"),
  2313 => (x"da",x"c2",x"87",x"c2"),
  2314 => (x"c1",x"4a",x"bf",x"cc"),
  2315 => (x"d0",x"da",x"c2",x"ba"),
  2316 => (x"7a",x"0a",x"fc",x"5a"),
  2317 => (x"c1",x"9a",x"c1",x"0a"),
  2318 => (x"e9",x"49",x"a2",x"c0"),
  2319 => (x"da",x"c1",x"87",x"da"),
  2320 => (x"87",x"e3",x"e6",x"49"),
  2321 => (x"da",x"c2",x"7e",x"c1"),
  2322 => (x"66",x"c8",x"48",x"c4"),
  2323 => (x"cc",x"da",x"c2",x"78"),
  2324 => (x"e9",x"c0",x"05",x"bf"),
  2325 => (x"c3",x"49",x"75",x"87"),
  2326 => (x"1e",x"71",x"99",x"ff"),
  2327 => (x"f8",x"fb",x"49",x"c0"),
  2328 => (x"c8",x"49",x"75",x"87"),
  2329 => (x"1e",x"71",x"29",x"b7"),
  2330 => (x"ec",x"fb",x"49",x"c1"),
  2331 => (x"c3",x"86",x"c8",x"87"),
  2332 => (x"f2",x"e5",x"49",x"fd"),
  2333 => (x"49",x"fa",x"c3",x"87"),
  2334 => (x"c7",x"87",x"ec",x"e5"),
  2335 => (x"49",x"75",x"87",x"f4"),
  2336 => (x"c8",x"99",x"ff",x"c3"),
  2337 => (x"b5",x"71",x"2d",x"b7"),
  2338 => (x"c0",x"02",x"9d",x"75"),
  2339 => (x"a6",x"c8",x"87",x"e4"),
  2340 => (x"bf",x"c8",x"ff",x"48"),
  2341 => (x"49",x"66",x"c8",x"78"),
  2342 => (x"bf",x"c8",x"da",x"c2"),
  2343 => (x"a9",x"e0",x"c2",x"89"),
  2344 => (x"87",x"c4",x"c0",x"03"),
  2345 => (x"87",x"d0",x"4d",x"c0"),
  2346 => (x"48",x"c8",x"da",x"c2"),
  2347 => (x"c0",x"78",x"66",x"c8"),
  2348 => (x"da",x"c2",x"87",x"c6"),
  2349 => (x"78",x"c0",x"48",x"c8"),
  2350 => (x"99",x"c8",x"49",x"75"),
  2351 => (x"87",x"ce",x"c0",x"05"),
  2352 => (x"e4",x"49",x"f5",x"c3"),
  2353 => (x"49",x"70",x"87",x"e1"),
  2354 => (x"c0",x"02",x"99",x"c2"),
  2355 => (x"ca",x"c3",x"87",x"e7"),
  2356 => (x"c0",x"02",x"bf",x"c4"),
  2357 => (x"c1",x"48",x"87",x"ca"),
  2358 => (x"c8",x"ca",x"c3",x"88"),
  2359 => (x"87",x"d3",x"c0",x"58"),
  2360 => (x"c1",x"48",x"66",x"c4"),
  2361 => (x"7e",x"70",x"80",x"e0"),
  2362 => (x"c0",x"02",x"bf",x"6e"),
  2363 => (x"ff",x"4b",x"87",x"c5"),
  2364 => (x"c1",x"0f",x"73",x"49"),
  2365 => (x"c4",x"49",x"75",x"7e"),
  2366 => (x"ce",x"c0",x"05",x"99"),
  2367 => (x"49",x"f2",x"c3",x"87"),
  2368 => (x"70",x"87",x"e4",x"e3"),
  2369 => (x"02",x"99",x"c2",x"49"),
  2370 => (x"c3",x"87",x"ea",x"c0"),
  2371 => (x"7e",x"bf",x"c4",x"ca"),
  2372 => (x"a8",x"b7",x"c7",x"48"),
  2373 => (x"87",x"cb",x"c0",x"03"),
  2374 => (x"80",x"c1",x"48",x"6e"),
  2375 => (x"58",x"c8",x"ca",x"c3"),
  2376 => (x"c4",x"87",x"d0",x"c0"),
  2377 => (x"e0",x"c1",x"4a",x"66"),
  2378 => (x"c0",x"02",x"6a",x"82"),
  2379 => (x"fe",x"4b",x"87",x"c5"),
  2380 => (x"c1",x"0f",x"73",x"49"),
  2381 => (x"49",x"fd",x"c3",x"7e"),
  2382 => (x"70",x"87",x"ec",x"e2"),
  2383 => (x"02",x"99",x"c2",x"49"),
  2384 => (x"c3",x"87",x"e6",x"c0"),
  2385 => (x"02",x"bf",x"c4",x"ca"),
  2386 => (x"c3",x"87",x"c9",x"c0"),
  2387 => (x"c0",x"48",x"c4",x"ca"),
  2388 => (x"87",x"d3",x"c0",x"78"),
  2389 => (x"c1",x"48",x"66",x"c4"),
  2390 => (x"7e",x"70",x"80",x"e0"),
  2391 => (x"c0",x"02",x"bf",x"6e"),
  2392 => (x"fd",x"4b",x"87",x"c5"),
  2393 => (x"c1",x"0f",x"73",x"49"),
  2394 => (x"49",x"fa",x"c3",x"7e"),
  2395 => (x"70",x"87",x"f8",x"e1"),
  2396 => (x"02",x"99",x"c2",x"49"),
  2397 => (x"c3",x"87",x"ea",x"c0"),
  2398 => (x"48",x"bf",x"c4",x"ca"),
  2399 => (x"03",x"a8",x"b7",x"c7"),
  2400 => (x"c3",x"87",x"c9",x"c0"),
  2401 => (x"c7",x"48",x"c4",x"ca"),
  2402 => (x"87",x"d3",x"c0",x"78"),
  2403 => (x"c1",x"48",x"66",x"c4"),
  2404 => (x"7e",x"70",x"80",x"e0"),
  2405 => (x"c0",x"02",x"bf",x"6e"),
  2406 => (x"fc",x"4b",x"87",x"c5"),
  2407 => (x"c1",x"0f",x"73",x"49"),
  2408 => (x"c3",x"48",x"75",x"7e"),
  2409 => (x"a6",x"cc",x"98",x"f0"),
  2410 => (x"05",x"98",x"70",x"58"),
  2411 => (x"c1",x"87",x"ce",x"c0"),
  2412 => (x"f2",x"e0",x"49",x"da"),
  2413 => (x"c2",x"49",x"70",x"87"),
  2414 => (x"f9",x"c1",x"02",x"99"),
  2415 => (x"49",x"e8",x"cf",x"87"),
  2416 => (x"70",x"87",x"cd",x"c3"),
  2417 => (x"fc",x"c9",x"c3",x"4b"),
  2418 => (x"c3",x"50",x"c0",x"48"),
  2419 => (x"bf",x"97",x"fc",x"c9"),
  2420 => (x"87",x"d2",x"c1",x"05"),
  2421 => (x"c0",x"05",x"66",x"c8"),
  2422 => (x"da",x"c1",x"87",x"cc"),
  2423 => (x"87",x"c7",x"e0",x"49"),
  2424 => (x"c1",x"02",x"98",x"70"),
  2425 => (x"bf",x"e8",x"87",x"c0"),
  2426 => (x"ff",x"c3",x"49",x"4d"),
  2427 => (x"2d",x"b7",x"c8",x"99"),
  2428 => (x"db",x"ff",x"b5",x"71"),
  2429 => (x"49",x"73",x"87",x"ea"),
  2430 => (x"70",x"87",x"e1",x"c2"),
  2431 => (x"c6",x"c0",x"02",x"98"),
  2432 => (x"fc",x"c9",x"c3",x"87"),
  2433 => (x"c3",x"50",x"c1",x"48"),
  2434 => (x"bf",x"97",x"fc",x"c9"),
  2435 => (x"87",x"d6",x"c0",x"05"),
  2436 => (x"f0",x"c3",x"49",x"75"),
  2437 => (x"cd",x"ff",x"05",x"99"),
  2438 => (x"49",x"da",x"c1",x"87"),
  2439 => (x"87",x"c7",x"df",x"ff"),
  2440 => (x"ff",x"05",x"98",x"70"),
  2441 => (x"ca",x"c3",x"87",x"c0"),
  2442 => (x"4b",x"49",x"bf",x"c4"),
  2443 => (x"66",x"c4",x"93",x"cc"),
  2444 => (x"71",x"4b",x"6b",x"83"),
  2445 => (x"9c",x"74",x"0f",x"73"),
  2446 => (x"87",x"e9",x"c0",x"02"),
  2447 => (x"e4",x"c0",x"02",x"6c"),
  2448 => (x"ff",x"49",x"6c",x"87"),
  2449 => (x"70",x"87",x"e0",x"de"),
  2450 => (x"02",x"99",x"c1",x"49"),
  2451 => (x"c4",x"87",x"cb",x"c0"),
  2452 => (x"ca",x"c3",x"4b",x"a4"),
  2453 => (x"6b",x"49",x"bf",x"c4"),
  2454 => (x"84",x"c8",x"0f",x"4b"),
  2455 => (x"87",x"c5",x"c0",x"02"),
  2456 => (x"dc",x"ff",x"05",x"6c"),
  2457 => (x"c0",x"02",x"6e",x"87"),
  2458 => (x"ca",x"c3",x"87",x"c8"),
  2459 => (x"f1",x"49",x"bf",x"c4"),
  2460 => (x"8e",x"f4",x"87",x"ea"),
  2461 => (x"4c",x"26",x"4d",x"26"),
  2462 => (x"4f",x"26",x"4b",x"26"),
  2463 => (x"00",x"00",x"00",x"10"),
  2464 => (x"00",x"00",x"00",x"00"),
  2465 => (x"00",x"00",x"00",x"00"),
  2466 => (x"00",x"00",x"00",x"00"),
  2467 => (x"00",x"00",x"00",x"00"),
  2468 => (x"ff",x"4a",x"71",x"1e"),
  2469 => (x"72",x"49",x"bf",x"c8"),
  2470 => (x"4f",x"26",x"48",x"a1"),
  2471 => (x"bf",x"c8",x"ff",x"1e"),
  2472 => (x"c0",x"c0",x"fe",x"89"),
  2473 => (x"a9",x"c0",x"c0",x"c0"),
  2474 => (x"c0",x"87",x"c4",x"01"),
  2475 => (x"c1",x"87",x"c2",x"4a"),
  2476 => (x"26",x"48",x"72",x"4a"),
  2477 => (x"5b",x"5e",x"0e",x"4f"),
  2478 => (x"71",x"0e",x"5d",x"5c"),
  2479 => (x"4c",x"d4",x"ff",x"4b"),
  2480 => (x"c0",x"48",x"66",x"d0"),
  2481 => (x"ff",x"49",x"d6",x"78"),
  2482 => (x"c3",x"87",x"d9",x"dd"),
  2483 => (x"49",x"6c",x"7c",x"ff"),
  2484 => (x"71",x"99",x"ff",x"c3"),
  2485 => (x"f0",x"c3",x"49",x"4d"),
  2486 => (x"a9",x"e0",x"c1",x"99"),
  2487 => (x"c3",x"87",x"cb",x"05"),
  2488 => (x"48",x"6c",x"7c",x"ff"),
  2489 => (x"66",x"d0",x"98",x"c3"),
  2490 => (x"ff",x"c3",x"78",x"08"),
  2491 => (x"49",x"4a",x"6c",x"7c"),
  2492 => (x"ff",x"c3",x"31",x"c8"),
  2493 => (x"71",x"4a",x"6c",x"7c"),
  2494 => (x"c8",x"49",x"72",x"b2"),
  2495 => (x"7c",x"ff",x"c3",x"31"),
  2496 => (x"b2",x"71",x"4a",x"6c"),
  2497 => (x"31",x"c8",x"49",x"72"),
  2498 => (x"6c",x"7c",x"ff",x"c3"),
  2499 => (x"ff",x"b2",x"71",x"4a"),
  2500 => (x"e0",x"c0",x"48",x"d0"),
  2501 => (x"02",x"9b",x"73",x"78"),
  2502 => (x"7b",x"72",x"87",x"c2"),
  2503 => (x"4d",x"26",x"48",x"75"),
  2504 => (x"4b",x"26",x"4c",x"26"),
  2505 => (x"26",x"1e",x"4f",x"26"),
  2506 => (x"5b",x"5e",x"0e",x"4f"),
  2507 => (x"86",x"f8",x"0e",x"5c"),
  2508 => (x"a6",x"c8",x"1e",x"76"),
  2509 => (x"87",x"fd",x"fd",x"49"),
  2510 => (x"4b",x"70",x"86",x"c4"),
  2511 => (x"a8",x"c2",x"48",x"6e"),
  2512 => (x"87",x"fb",x"c2",x"03"),
  2513 => (x"f0",x"c3",x"4a",x"73"),
  2514 => (x"aa",x"d0",x"c1",x"9a"),
  2515 => (x"c1",x"87",x"c7",x"02"),
  2516 => (x"c2",x"05",x"aa",x"e0"),
  2517 => (x"49",x"73",x"87",x"e9"),
  2518 => (x"c3",x"02",x"99",x"c8"),
  2519 => (x"87",x"c6",x"ff",x"87"),
  2520 => (x"9c",x"c3",x"4c",x"73"),
  2521 => (x"c1",x"05",x"ac",x"c2"),
  2522 => (x"66",x"c4",x"87",x"c4"),
  2523 => (x"71",x"31",x"c9",x"49"),
  2524 => (x"4a",x"66",x"c4",x"1e"),
  2525 => (x"c3",x"92",x"cc",x"c1"),
  2526 => (x"72",x"49",x"cc",x"ca"),
  2527 => (x"cb",x"cd",x"fe",x"81"),
  2528 => (x"ff",x"49",x"d8",x"87"),
  2529 => (x"c8",x"87",x"dd",x"da"),
  2530 => (x"f6",x"c2",x"1e",x"c0"),
  2531 => (x"e6",x"fd",x"49",x"e8"),
  2532 => (x"d0",x"ff",x"87",x"e1"),
  2533 => (x"78",x"e0",x"c0",x"48"),
  2534 => (x"1e",x"e8",x"f6",x"c2"),
  2535 => (x"c1",x"4a",x"66",x"cc"),
  2536 => (x"ca",x"c3",x"92",x"cc"),
  2537 => (x"81",x"72",x"49",x"cc"),
  2538 => (x"87",x"e1",x"cb",x"fe"),
  2539 => (x"ac",x"c1",x"86",x"cc"),
  2540 => (x"87",x"cb",x"c1",x"05"),
  2541 => (x"fd",x"49",x"ee",x"c0"),
  2542 => (x"c4",x"87",x"d1",x"e3"),
  2543 => (x"31",x"c9",x"49",x"66"),
  2544 => (x"66",x"c4",x"1e",x"71"),
  2545 => (x"92",x"cc",x"c1",x"4a"),
  2546 => (x"49",x"cc",x"ca",x"c3"),
  2547 => (x"cb",x"fe",x"81",x"72"),
  2548 => (x"f6",x"c2",x"87",x"fa"),
  2549 => (x"66",x"c8",x"1e",x"e8"),
  2550 => (x"92",x"cc",x"c1",x"4a"),
  2551 => (x"49",x"cc",x"ca",x"c3"),
  2552 => (x"c9",x"fe",x"81",x"72"),
  2553 => (x"49",x"d7",x"87",x"e8"),
  2554 => (x"87",x"f8",x"d8",x"ff"),
  2555 => (x"c2",x"1e",x"c0",x"c8"),
  2556 => (x"fd",x"49",x"e8",x"f6"),
  2557 => (x"cc",x"87",x"d9",x"e4"),
  2558 => (x"48",x"d0",x"ff",x"86"),
  2559 => (x"f8",x"78",x"e0",x"c0"),
  2560 => (x"26",x"4c",x"26",x"8e"),
  2561 => (x"1e",x"4f",x"26",x"4b"),
  2562 => (x"b7",x"c2",x"4a",x"71"),
  2563 => (x"87",x"ce",x"03",x"aa"),
  2564 => (x"cc",x"c1",x"49",x"72"),
  2565 => (x"cc",x"ca",x"c3",x"91"),
  2566 => (x"81",x"c8",x"c1",x"81"),
  2567 => (x"4f",x"26",x"79",x"c0"),
  2568 => (x"5c",x"5b",x"5e",x"0e"),
  2569 => (x"86",x"fc",x"0e",x"5d"),
  2570 => (x"d4",x"ff",x"4a",x"71"),
  2571 => (x"d4",x"4c",x"c0",x"4b"),
  2572 => (x"b7",x"c3",x"4d",x"66"),
  2573 => (x"c2",x"c2",x"01",x"ad"),
  2574 => (x"02",x"9a",x"72",x"87"),
  2575 => (x"1e",x"87",x"ec",x"c0"),
  2576 => (x"cc",x"c1",x"49",x"75"),
  2577 => (x"cc",x"ca",x"c3",x"91"),
  2578 => (x"c8",x"80",x"71",x"48"),
  2579 => (x"66",x"c4",x"58",x"a6"),
  2580 => (x"c3",x"c3",x"fe",x"49"),
  2581 => (x"70",x"86",x"c4",x"87"),
  2582 => (x"87",x"d4",x"02",x"98"),
  2583 => (x"c8",x"c1",x"49",x"6e"),
  2584 => (x"6e",x"79",x"c1",x"81"),
  2585 => (x"69",x"81",x"c8",x"49"),
  2586 => (x"75",x"87",x"c5",x"4c"),
  2587 => (x"87",x"d7",x"fe",x"49"),
  2588 => (x"c8",x"48",x"d0",x"ff"),
  2589 => (x"7b",x"dd",x"78",x"e1"),
  2590 => (x"ff",x"c3",x"48",x"74"),
  2591 => (x"74",x"7b",x"70",x"98"),
  2592 => (x"29",x"b7",x"c8",x"49"),
  2593 => (x"ff",x"c3",x"48",x"71"),
  2594 => (x"74",x"7b",x"70",x"98"),
  2595 => (x"29",x"b7",x"d0",x"49"),
  2596 => (x"ff",x"c3",x"48",x"71"),
  2597 => (x"74",x"7b",x"70",x"98"),
  2598 => (x"28",x"b7",x"d8",x"48"),
  2599 => (x"7b",x"c0",x"7b",x"70"),
  2600 => (x"7b",x"7b",x"7b",x"7b"),
  2601 => (x"7b",x"7b",x"7b",x"7b"),
  2602 => (x"ff",x"7b",x"7b",x"7b"),
  2603 => (x"e0",x"c0",x"48",x"d0"),
  2604 => (x"dc",x"1e",x"75",x"78"),
  2605 => (x"d0",x"d6",x"ff",x"49"),
  2606 => (x"fc",x"86",x"c4",x"87"),
  2607 => (x"26",x"4d",x"26",x"8e"),
  2608 => (x"26",x"4b",x"26",x"4c"),
  2609 => (x"d4",x"ff",x"1e",x"4f"),
  2610 => (x"7a",x"ff",x"c3",x"4a"),
  2611 => (x"c5",x"48",x"d0",x"ff"),
  2612 => (x"71",x"7a",x"c4",x"78"),
  2613 => (x"28",x"b7",x"d8",x"48"),
  2614 => (x"48",x"71",x"7a",x"70"),
  2615 => (x"70",x"28",x"b7",x"d0"),
  2616 => (x"c8",x"48",x"71",x"7a"),
  2617 => (x"7a",x"70",x"28",x"b7"),
  2618 => (x"d0",x"ff",x"7a",x"71"),
  2619 => (x"26",x"78",x"c4",x"48"),
  2620 => (x"4a",x"c0",x"1e",x"4f"),
  2621 => (x"bf",x"e4",x"cc",x"c3"),
  2622 => (x"49",x"87",x"ca",x"02"),
  2623 => (x"48",x"e4",x"cc",x"c3"),
  2624 => (x"11",x"78",x"a1",x"c1"),
  2625 => (x"05",x"9a",x"72",x"4a"),
  2626 => (x"cc",x"c3",x"87",x"c6"),
  2627 => (x"78",x"c0",x"48",x"e4"),
  2628 => (x"4f",x"26",x"48",x"72"),
  2629 => (x"e4",x"cc",x"c3",x"1e"),
  2630 => (x"c0",x"eb",x"c2",x"48"),
  2631 => (x"4f",x"26",x"78",x"bf"),
  2632 => (x"5c",x"5b",x"5e",x"0e"),
  2633 => (x"ff",x"4a",x"71",x"0e"),
  2634 => (x"d4",x"ff",x"4c",x"d0"),
  2635 => (x"c1",x"7c",x"c5",x"4b"),
  2636 => (x"7b",x"c3",x"7b",x"d5"),
  2637 => (x"7c",x"c5",x"7c",x"c4"),
  2638 => (x"c1",x"7b",x"d3",x"c1"),
  2639 => (x"c8",x"7c",x"c4",x"7b"),
  2640 => (x"d4",x"c1",x"7c",x"c5"),
  2641 => (x"b7",x"49",x"c0",x"7b"),
  2642 => (x"87",x"ca",x"06",x"aa"),
  2643 => (x"81",x"c1",x"7b",x"c0"),
  2644 => (x"04",x"a9",x"b7",x"72"),
  2645 => (x"7c",x"c4",x"87",x"f6"),
  2646 => (x"d3",x"c1",x"7c",x"c5"),
  2647 => (x"c4",x"7b",x"c0",x"7b"),
  2648 => (x"26",x"4c",x"26",x"7c"),
  2649 => (x"1e",x"4f",x"26",x"4b"),
  2650 => (x"4b",x"71",x"1e",x"73"),
  2651 => (x"fc",x"c3",x"c3",x"1e"),
  2652 => (x"e3",x"fe",x"fd",x"49"),
  2653 => (x"70",x"86",x"c4",x"87"),
  2654 => (x"e1",x"c0",x"02",x"98"),
  2655 => (x"c4",x"c4",x"c3",x"87"),
  2656 => (x"2a",x"ca",x"4a",x"bf"),
  2657 => (x"02",x"8a",x"c0",x"c3"),
  2658 => (x"c0",x"c1",x"87",x"ce"),
  2659 => (x"87",x"ce",x"05",x"8a"),
  2660 => (x"48",x"dc",x"e8",x"c1"),
  2661 => (x"87",x"c6",x"50",x"c0"),
  2662 => (x"48",x"dc",x"e8",x"c1"),
  2663 => (x"4b",x"26",x"50",x"c1"),
  2664 => (x"73",x"1e",x"4f",x"26"),
  2665 => (x"f8",x"c3",x"c3",x"1e"),
  2666 => (x"c1",x"50",x"c0",x"48"),
  2667 => (x"c1",x"48",x"dc",x"e8"),
  2668 => (x"c4",x"ff",x"c0",x"50"),
  2669 => (x"c1",x"50",x"c0",x"48"),
  2670 => (x"87",x"c9",x"fc",x"49"),
  2671 => (x"49",x"c0",x"c0",x"c4"),
  2672 => (x"c2",x"87",x"dd",x"fd"),
  2673 => (x"49",x"bf",x"d4",x"eb"),
  2674 => (x"c2",x"87",x"dc",x"fe"),
  2675 => (x"49",x"bf",x"d4",x"eb"),
  2676 => (x"87",x"d6",x"d8",x"fe"),
  2677 => (x"ec",x"fb",x"49",x"c0"),
  2678 => (x"49",x"d0",x"c6",x"87"),
  2679 => (x"70",x"87",x"f1",x"f2"),
  2680 => (x"f7",x"f2",x"49",x"4b"),
  2681 => (x"05",x"98",x"70",x"87"),
  2682 => (x"49",x"73",x"87",x"ca"),
  2683 => (x"70",x"87",x"ed",x"f2"),
  2684 => (x"87",x"f6",x"02",x"98"),
  2685 => (x"cc",x"fb",x"49",x"c1"),
  2686 => (x"49",x"e4",x"c1",x"87"),
  2687 => (x"70",x"87",x"d1",x"f2"),
  2688 => (x"d7",x"f2",x"49",x"4b"),
  2689 => (x"05",x"98",x"70",x"87"),
  2690 => (x"49",x"73",x"87",x"ca"),
  2691 => (x"70",x"87",x"cd",x"f2"),
  2692 => (x"87",x"f6",x"02",x"98"),
  2693 => (x"ec",x"fa",x"49",x"c0"),
  2694 => (x"26",x"48",x"c0",x"87"),
  2695 => (x"1e",x"4f",x"26",x"4b"),
  2696 => (x"ea",x"c2",x"1e",x"73"),
  2697 => (x"c0",x"05",x"bf",x"fc"),
  2698 => (x"c9",x"c3",x"87",x"ea"),
  2699 => (x"c4",x"ff",x"49",x"d8"),
  2700 => (x"b7",x"c0",x"87",x"e8"),
  2701 => (x"87",x"ce",x"04",x"a8"),
  2702 => (x"49",x"d8",x"c9",x"c3"),
  2703 => (x"87",x"da",x"c4",x"ff"),
  2704 => (x"03",x"a8",x"b7",x"c0"),
  2705 => (x"ea",x"c2",x"87",x"f2"),
  2706 => (x"c1",x"48",x"bf",x"fc"),
  2707 => (x"c0",x"eb",x"c2",x"80"),
  2708 => (x"87",x"e2",x"c1",x"58"),
  2709 => (x"bf",x"fc",x"ea",x"c2"),
  2710 => (x"99",x"c1",x"49",x"4b"),
  2711 => (x"87",x"f0",x"c0",x"02"),
  2712 => (x"b7",x"c1",x"49",x"73"),
  2713 => (x"d8",x"eb",x"c2",x"29"),
  2714 => (x"9a",x"4a",x"11",x"81"),
  2715 => (x"87",x"c6",x"c1",x"02"),
  2716 => (x"06",x"aa",x"b7",x"c1"),
  2717 => (x"1e",x"72",x"87",x"cc"),
  2718 => (x"49",x"d8",x"c9",x"c3"),
  2719 => (x"87",x"e6",x"c1",x"ff"),
  2720 => (x"ea",x"c2",x"86",x"c4"),
  2721 => (x"c1",x"48",x"bf",x"fc"),
  2722 => (x"c0",x"eb",x"c2",x"80"),
  2723 => (x"87",x"e6",x"c0",x"58"),
  2724 => (x"49",x"d8",x"c9",x"c3"),
  2725 => (x"87",x"c2",x"c3",x"ff"),
  2726 => (x"ea",x"c2",x"4a",x"70"),
  2727 => (x"87",x"cb",x"02",x"aa"),
  2728 => (x"02",x"aa",x"fa",x"c3"),
  2729 => (x"aa",x"c3",x"87",x"c5"),
  2730 => (x"c2",x"87",x"cb",x"05"),
  2731 => (x"48",x"bf",x"fc",x"ea"),
  2732 => (x"eb",x"c2",x"80",x"c1"),
  2733 => (x"4b",x"26",x"58",x"c0"),
  2734 => (x"00",x"00",x"4f",x"26"),
  2735 => (x"00",x"00",x"00",x"00"),
  2736 => (x"00",x"00",x"2b",x"f0"),
  2737 => (x"11",x"14",x"12",x"58"),
  2738 => (x"23",x"1c",x"1b",x"1d"),
  2739 => (x"91",x"94",x"59",x"5a"),
  2740 => (x"f4",x"eb",x"f2",x"f5"),
  2741 => (x"00",x"00",x"2d",x"68"),
  2742 => (x"f3",x"c8",x"f3",x"ff"),
  2743 => (x"f2",x"50",x"f3",x"64"),
  2744 => (x"1e",x"00",x"f4",x"01"),
  2745 => (x"4b",x"71",x"1e",x"73"),
  2746 => (x"c5",x"e8",x"fe",x"49"),
  2747 => (x"fc",x"c9",x"c3",x"87"),
  2748 => (x"c7",x"02",x"bf",x"97"),
  2749 => (x"c0",x"c0",x"c4",x"87"),
  2750 => (x"87",x"e4",x"f8",x"49"),
  2751 => (x"e7",x"fe",x"49",x"73"),
  2752 => (x"4b",x"26",x"87",x"f0"),
  2753 => (x"73",x"1e",x"4f",x"26"),
  2754 => (x"c3",x"4a",x"71",x"1e"),
  2755 => (x"4b",x"bf",x"f0",x"c3"),
  2756 => (x"c5",x"02",x"9a",x"72"),
  2757 => (x"bb",x"c0",x"c2",x"87"),
  2758 => (x"c0",x"c1",x"87",x"c3"),
  2759 => (x"f6",x"49",x"73",x"bb"),
  2760 => (x"f4",x"c7",x"87",x"e3"),
  2761 => (x"87",x"e8",x"ed",x"49"),
  2762 => (x"ed",x"49",x"4b",x"70"),
  2763 => (x"98",x"70",x"87",x"ee"),
  2764 => (x"73",x"87",x"ca",x"05"),
  2765 => (x"87",x"e4",x"ed",x"49"),
  2766 => (x"f6",x"02",x"98",x"70"),
  2767 => (x"26",x"4b",x"26",x"87"),
  2768 => (x"5b",x"5e",x"0e",x"4f"),
  2769 => (x"4b",x"71",x"0e",x"5c"),
  2770 => (x"d3",x"02",x"66",x"cc"),
  2771 => (x"f0",x"c0",x"4c",x"87"),
  2772 => (x"e9",x"c0",x"02",x"8c"),
  2773 => (x"c1",x"49",x"74",x"87"),
  2774 => (x"e1",x"c0",x"02",x"89"),
  2775 => (x"87",x"f3",x"c0",x"87"),
  2776 => (x"c0",x"02",x"9b",x"73"),
  2777 => (x"c3",x"c3",x"87",x"ed"),
  2778 => (x"c1",x"49",x"bf",x"f0"),
  2779 => (x"d4",x"f5",x"71",x"b1"),
  2780 => (x"f7",x"49",x"73",x"87"),
  2781 => (x"49",x"73",x"87",x"f1"),
  2782 => (x"87",x"ee",x"d1",x"fe"),
  2783 => (x"1e",x"74",x"87",x"d5"),
  2784 => (x"db",x"f2",x"49",x"c0"),
  2785 => (x"fd",x"49",x"74",x"87"),
  2786 => (x"1e",x"74",x"87",x"fc"),
  2787 => (x"cf",x"f2",x"49",x"73"),
  2788 => (x"c3",x"86",x"c8",x"87"),
  2789 => (x"49",x"bf",x"f0",x"c3"),
  2790 => (x"26",x"87",x"ea",x"f4"),
  2791 => (x"26",x"4b",x"26",x"4c"),
  2792 => (x"c4",x"ff",x"1e",x"4f"),
  2793 => (x"d4",x"ff",x"87",x"df"),
  2794 => (x"78",x"ff",x"c3",x"48"),
  2795 => (x"87",x"d0",x"df",x"fd"),
  2796 => (x"cd",x"02",x"98",x"70"),
  2797 => (x"ee",x"e8",x"fd",x"87"),
  2798 => (x"02",x"98",x"70",x"87"),
  2799 => (x"4a",x"c1",x"87",x"c4"),
  2800 => (x"4a",x"c0",x"87",x"c2"),
  2801 => (x"c8",x"02",x"9a",x"72"),
  2802 => (x"ec",x"ef",x"c2",x"87"),
  2803 => (x"d6",x"d3",x"fd",x"49"),
  2804 => (x"fe",x"49",x"c0",x"87"),
  2805 => (x"f7",x"87",x"e1",x"f8"),
  2806 => (x"fb",x"fe",x"87",x"c8"),
  2807 => (x"fe",x"f8",x"87",x"e1"),
  2808 => (x"e5",x"de",x"ff",x"87"),
  2809 => (x"87",x"c1",x"ed",x"87"),
  2810 => (x"4f",x"26",x"87",x"f4"),
  2811 => (x"00",x"00",x"4b",x"4f"),
  2812 => (x"72",x"61",x"74",x"41"),
  2813 => (x"54",x"53",x"20",x"69"),
  2814 => (x"30",x"53",x"3b",x"3b"),
  2815 => (x"54",x"53",x"2c",x"55"),
  2816 => (x"6c",x"46",x"2c",x"20"),
  2817 => (x"79",x"70",x"70",x"6f"),
  2818 => (x"3b",x"3a",x"41",x"20"),
  2819 => (x"2c",x"55",x"31",x"53"),
  2820 => (x"2c",x"20",x"54",x"53"),
  2821 => (x"70",x"6f",x"6c",x"46"),
  2822 => (x"42",x"20",x"79",x"70"),
  2823 => (x"36",x"4f",x"3b",x"3a"),
  2824 => (x"72",x"57",x"2c",x"37"),
  2825 => (x"20",x"65",x"74",x"69"),
  2826 => (x"74",x"6f",x"72",x"70"),
  2827 => (x"2c",x"74",x"63",x"65"),
  2828 => (x"2c",x"66",x"66",x"4f"),
  2829 => (x"42",x"2c",x"3a",x"41"),
  2830 => (x"6f",x"42",x"2c",x"3a"),
  2831 => (x"46",x"3b",x"68",x"74"),
  2832 => (x"47",x"4d",x"49",x"2c"),
  2833 => (x"2c",x"4d",x"4f",x"52"),
  2834 => (x"64",x"61",x"6f",x"4c"),
  2835 => (x"4d",x"4f",x"52",x"20"),
  2836 => (x"2c",x"31",x"50",x"3b"),
  2837 => (x"43",x"20",x"54",x"53"),
  2838 => (x"69",x"66",x"6e",x"6f"),
  2839 => (x"61",x"72",x"75",x"67"),
  2840 => (x"6e",x"6f",x"69",x"74"),
  2841 => (x"4f",x"31",x"50",x"3b"),
  2842 => (x"52",x"2c",x"33",x"31"),
  2843 => (x"28",x"20",x"4d",x"41"),
  2844 => (x"64",x"65",x"65",x"6e"),
  2845 => (x"72",x"61",x"48",x"20"),
  2846 => (x"65",x"52",x"20",x"64"),
  2847 => (x"29",x"74",x"65",x"73"),
  2848 => (x"32",x"31",x"35",x"2c"),
  2849 => (x"4d",x"31",x"2c",x"4b"),
  2850 => (x"4d",x"32",x"2c",x"42"),
  2851 => (x"4d",x"34",x"2c",x"42"),
  2852 => (x"4d",x"38",x"2c",x"42"),
  2853 => (x"34",x"31",x"2c",x"42"),
  2854 => (x"50",x"3b",x"42",x"4d"),
  2855 => (x"2c",x"38",x"4f",x"31"),
  2856 => (x"65",x"64",x"69",x"56"),
  2857 => (x"6f",x"6d",x"20",x"6f"),
  2858 => (x"4d",x"2c",x"65",x"64"),
  2859 => (x"2c",x"6f",x"6e",x"6f"),
  2860 => (x"6f",x"6c",x"6f",x"43"),
  2861 => (x"50",x"3b",x"72",x"75"),
  2862 => (x"4f",x"4e",x"4f",x"31"),
  2863 => (x"69",x"68",x"43",x"2c"),
  2864 => (x"74",x"65",x"73",x"70"),
  2865 => (x"2c",x"54",x"53",x"2c"),
  2866 => (x"2c",x"45",x"54",x"53"),
  2867 => (x"61",x"67",x"65",x"4d"),
  2868 => (x"3b",x"45",x"54",x"53"),
  2869 => (x"4a",x"4f",x"31",x"50"),
  2870 => (x"20",x"54",x"53",x"2c"),
  2871 => (x"74",x"69",x"6c",x"42"),
  2872 => (x"2c",x"72",x"65",x"74"),
  2873 => (x"2c",x"66",x"66",x"4f"),
  2874 => (x"50",x"3b",x"6e",x"4f"),
  2875 => (x"2c",x"4d",x"4f",x"31"),
  2876 => (x"72",x"65",x"74",x"53"),
  2877 => (x"73",x"20",x"6f",x"65"),
  2878 => (x"64",x"6e",x"75",x"6f"),
  2879 => (x"66",x"66",x"4f",x"2c"),
  2880 => (x"3b",x"6e",x"4f",x"2c"),
  2881 => (x"4b",x"4f",x"31",x"50"),
  2882 => (x"63",x"53",x"2c",x"4c"),
  2883 => (x"69",x"6c",x"6e",x"61"),
  2884 => (x"2c",x"73",x"65",x"6e"),
  2885 => (x"2c",x"66",x"66",x"4f"),
  2886 => (x"2c",x"25",x"35",x"32"),
  2887 => (x"2c",x"25",x"30",x"35"),
  2888 => (x"3b",x"25",x"35",x"37"),
  2889 => (x"54",x"4f",x"31",x"50"),
  2890 => (x"6d",x"6f",x"43",x"2c"),
  2891 => (x"69",x"73",x"6f",x"70"),
  2892 => (x"62",x"20",x"65",x"74"),
  2893 => (x"64",x"6e",x"65",x"6c"),
  2894 => (x"66",x"66",x"4f",x"2c"),
  2895 => (x"3b",x"6e",x"4f",x"2c"),
  2896 => (x"52",x"2c",x"30",x"54"),
  2897 => (x"74",x"65",x"73",x"65"),
  2898 => (x"6f",x"48",x"28",x"20"),
  2899 => (x"66",x"20",x"64",x"6c"),
  2900 => (x"68",x"20",x"72",x"6f"),
  2901 => (x"20",x"64",x"72",x"61"),
  2902 => (x"65",x"73",x"65",x"72"),
  2903 => (x"56",x"3b",x"29",x"74"),
  2904 => (x"2e",x"33",x"76",x"2c"),
  2905 => (x"00",x"2e",x"30",x"34"),
  2906 => (x"20",x"53",x"4f",x"54"),
  2907 => (x"20",x"20",x"20",x"20"),
  2908 => (x"00",x"47",x"4d",x"49"),
  2909 => (x"00",x"00",x"1a",x"af"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

